module network_tb;
 parameter DataSize=8'd172;
    parameter PayloadLen=128;
    parameter DataWidth=256;
    parameter WeightPos=144;
    parameter WeightWidth=8;
    parameter IndexPos=128;
    parameter IndexWidth=16;
    parameter PriorityPos=152;
    parameter PriorityWidth=8;
    parameter ExitPos=160;
    parameter ExitWidth=4;
    parameter InterNodeFIFODepth=256;
    parameter IntraNodeFIFODepth=1;
    parameter RoutingTableWidth=32;
    parameter RoutingTablesize=16;
    parameter MulticastTableWidth=103;
    parameter MulticastTablesize=16;
    parameter ReductionTableWidth=170;
    parameter ReductionTablesize=16;
    parameter PcktTypeLen=4;
    parameter LinkDelay=20;


 	reg clk,rst;

	always #5 clk=~clk;

	network#(
        .DataSize(DataSize),
        .PayloadLen(PayloadLen),
        .DataWidth(DataWidth),
        .WeightPos(WeightPos),
        .WeightWidth(WeightWidth),
        .IndexPos(IndexPos),
        .IndexWidth(IndexWidth),
        .PriorityPos(PriorityPos),
        .PriorityWidth(PriorityWidth),
        .ExitPos(ExitPos),
        .ExitWidth(ExitWidth),
        .InterNodeFIFODepth(InterNodeFIFODepth),
        .IntraNodeFIFODepth(IntraNodeFIFODepth),
        .RoutingTableWidth(RoutingTableWidth),
        .RoutingTablesize(RoutingTablesize),
        .MulticastTableWidth(MulticastTableWidth),
        .MulticastTablesize(MulticastTablesize),
        .ReductionTableWidth(ReductionTableWidth),
        .ReductionTablesize(ReductionTablesize),
        .PcktTypeLen(PcktTypeLen),
        .LinkDelay(LinkDelay)
    )
    net0(clk,rst);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_0_LOCAL.txt",net0.n_0_0_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_0_LOCAL.txt",net0.n_0_0_0.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_0_XPOS.txt",net0.n_0_0_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_0_XNEG.txt",net0.n_0_0_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_0_YPOS.txt",net0.n_0_0_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_0_YNEG.txt",net0.n_0_0_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_0_ZPOS.txt",net0.n_0_0_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_0_ZNEG.txt",net0.n_0_0_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_0_LOCAL.txt",net0.n_0_0_0.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_0_XPOS.txt",net0.n_0_0_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_0_XNEG.txt",net0.n_0_0_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_0_YPOS.txt",net0.n_0_0_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_0_YNEG.txt",net0.n_0_0_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_0_ZPOS.txt",net0.n_0_0_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_0_ZNEG.txt",net0.n_0_0_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_0_LOCAL.txt",net0.n_0_0_0.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_0_XPOS.txt",net0.n_0_0_0.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_0_XNEG.txt",net0.n_0_0_0.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_0_YPOS.txt",net0.n_0_0_0.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_0_YNEG.txt",net0.n_0_0_0.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_0_ZPOS.txt",net0.n_0_0_0.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_0_ZNEG.txt",net0.n_0_0_0.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_0_0_0.txt",net0.n_0_0_0.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_1_LOCAL.txt",net0.n_0_0_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_1_LOCAL.txt",net0.n_0_0_1.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_1_XPOS.txt",net0.n_0_0_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_1_XNEG.txt",net0.n_0_0_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_1_YPOS.txt",net0.n_0_0_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_1_YNEG.txt",net0.n_0_0_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_1_ZPOS.txt",net0.n_0_0_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_1_ZNEG.txt",net0.n_0_0_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_1_LOCAL.txt",net0.n_0_0_1.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_1_XPOS.txt",net0.n_0_0_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_1_XNEG.txt",net0.n_0_0_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_1_YPOS.txt",net0.n_0_0_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_1_YNEG.txt",net0.n_0_0_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_1_ZPOS.txt",net0.n_0_0_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_1_ZNEG.txt",net0.n_0_0_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_1_LOCAL.txt",net0.n_0_0_1.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_1_XPOS.txt",net0.n_0_0_1.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_1_XNEG.txt",net0.n_0_0_1.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_1_YPOS.txt",net0.n_0_0_1.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_1_YNEG.txt",net0.n_0_0_1.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_1_ZPOS.txt",net0.n_0_0_1.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_1_ZNEG.txt",net0.n_0_0_1.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_0_0_1.txt",net0.n_0_0_1.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_2_LOCAL.txt",net0.n_0_0_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_2_LOCAL.txt",net0.n_0_0_2.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_2_XPOS.txt",net0.n_0_0_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_2_XNEG.txt",net0.n_0_0_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_2_YPOS.txt",net0.n_0_0_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_2_YNEG.txt",net0.n_0_0_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_2_ZPOS.txt",net0.n_0_0_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_2_ZNEG.txt",net0.n_0_0_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_2_LOCAL.txt",net0.n_0_0_2.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_2_XPOS.txt",net0.n_0_0_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_2_XNEG.txt",net0.n_0_0_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_2_YPOS.txt",net0.n_0_0_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_2_YNEG.txt",net0.n_0_0_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_2_ZPOS.txt",net0.n_0_0_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_2_ZNEG.txt",net0.n_0_0_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_2_LOCAL.txt",net0.n_0_0_2.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_2_XPOS.txt",net0.n_0_0_2.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_2_XNEG.txt",net0.n_0_0_2.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_2_YPOS.txt",net0.n_0_0_2.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_2_YNEG.txt",net0.n_0_0_2.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_2_ZPOS.txt",net0.n_0_0_2.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_2_ZNEG.txt",net0.n_0_0_2.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_0_0_2.txt",net0.n_0_0_2.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_3_LOCAL.txt",net0.n_0_0_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_3_LOCAL.txt",net0.n_0_0_3.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_3_XPOS.txt",net0.n_0_0_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_3_XNEG.txt",net0.n_0_0_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_3_YPOS.txt",net0.n_0_0_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_3_YNEG.txt",net0.n_0_0_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_3_ZPOS.txt",net0.n_0_0_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_0_3_ZNEG.txt",net0.n_0_0_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_3_LOCAL.txt",net0.n_0_0_3.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_3_XPOS.txt",net0.n_0_0_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_3_XNEG.txt",net0.n_0_0_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_3_YPOS.txt",net0.n_0_0_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_3_YNEG.txt",net0.n_0_0_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_3_ZPOS.txt",net0.n_0_0_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_0_3_ZNEG.txt",net0.n_0_0_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_3_LOCAL.txt",net0.n_0_0_3.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_3_XPOS.txt",net0.n_0_0_3.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_3_XNEG.txt",net0.n_0_0_3.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_3_YPOS.txt",net0.n_0_0_3.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_3_YNEG.txt",net0.n_0_0_3.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_3_ZPOS.txt",net0.n_0_0_3.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_0_3_ZNEG.txt",net0.n_0_0_3.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_0_0_3.txt",net0.n_0_0_3.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_0_LOCAL.txt",net0.n_0_1_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_0_LOCAL.txt",net0.n_0_1_0.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_0_XPOS.txt",net0.n_0_1_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_0_XNEG.txt",net0.n_0_1_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_0_YPOS.txt",net0.n_0_1_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_0_YNEG.txt",net0.n_0_1_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_0_ZPOS.txt",net0.n_0_1_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_0_ZNEG.txt",net0.n_0_1_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_0_LOCAL.txt",net0.n_0_1_0.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_0_XPOS.txt",net0.n_0_1_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_0_XNEG.txt",net0.n_0_1_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_0_YPOS.txt",net0.n_0_1_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_0_YNEG.txt",net0.n_0_1_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_0_ZPOS.txt",net0.n_0_1_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_0_ZNEG.txt",net0.n_0_1_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_0_LOCAL.txt",net0.n_0_1_0.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_0_XPOS.txt",net0.n_0_1_0.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_0_XNEG.txt",net0.n_0_1_0.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_0_YPOS.txt",net0.n_0_1_0.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_0_YNEG.txt",net0.n_0_1_0.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_0_ZPOS.txt",net0.n_0_1_0.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_0_ZNEG.txt",net0.n_0_1_0.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_0_1_0.txt",net0.n_0_1_0.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_1_LOCAL.txt",net0.n_0_1_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_1_LOCAL.txt",net0.n_0_1_1.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_1_XPOS.txt",net0.n_0_1_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_1_XNEG.txt",net0.n_0_1_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_1_YPOS.txt",net0.n_0_1_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_1_YNEG.txt",net0.n_0_1_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_1_ZPOS.txt",net0.n_0_1_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_1_ZNEG.txt",net0.n_0_1_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_1_LOCAL.txt",net0.n_0_1_1.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_1_XPOS.txt",net0.n_0_1_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_1_XNEG.txt",net0.n_0_1_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_1_YPOS.txt",net0.n_0_1_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_1_YNEG.txt",net0.n_0_1_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_1_ZPOS.txt",net0.n_0_1_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_1_ZNEG.txt",net0.n_0_1_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_1_LOCAL.txt",net0.n_0_1_1.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_1_XPOS.txt",net0.n_0_1_1.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_1_XNEG.txt",net0.n_0_1_1.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_1_YPOS.txt",net0.n_0_1_1.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_1_YNEG.txt",net0.n_0_1_1.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_1_ZPOS.txt",net0.n_0_1_1.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_1_ZNEG.txt",net0.n_0_1_1.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_0_1_1.txt",net0.n_0_1_1.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_2_LOCAL.txt",net0.n_0_1_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_2_LOCAL.txt",net0.n_0_1_2.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_2_XPOS.txt",net0.n_0_1_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_2_XNEG.txt",net0.n_0_1_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_2_YPOS.txt",net0.n_0_1_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_2_YNEG.txt",net0.n_0_1_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_2_ZPOS.txt",net0.n_0_1_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_2_ZNEG.txt",net0.n_0_1_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_2_LOCAL.txt",net0.n_0_1_2.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_2_XPOS.txt",net0.n_0_1_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_2_XNEG.txt",net0.n_0_1_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_2_YPOS.txt",net0.n_0_1_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_2_YNEG.txt",net0.n_0_1_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_2_ZPOS.txt",net0.n_0_1_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_2_ZNEG.txt",net0.n_0_1_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_2_LOCAL.txt",net0.n_0_1_2.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_2_XPOS.txt",net0.n_0_1_2.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_2_XNEG.txt",net0.n_0_1_2.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_2_YPOS.txt",net0.n_0_1_2.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_2_YNEG.txt",net0.n_0_1_2.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_2_ZPOS.txt",net0.n_0_1_2.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_2_ZNEG.txt",net0.n_0_1_2.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_0_1_2.txt",net0.n_0_1_2.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_3_LOCAL.txt",net0.n_0_1_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_3_LOCAL.txt",net0.n_0_1_3.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_3_XPOS.txt",net0.n_0_1_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_3_XNEG.txt",net0.n_0_1_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_3_YPOS.txt",net0.n_0_1_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_3_YNEG.txt",net0.n_0_1_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_3_ZPOS.txt",net0.n_0_1_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_1_3_ZNEG.txt",net0.n_0_1_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_3_LOCAL.txt",net0.n_0_1_3.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_3_XPOS.txt",net0.n_0_1_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_3_XNEG.txt",net0.n_0_1_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_3_YPOS.txt",net0.n_0_1_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_3_YNEG.txt",net0.n_0_1_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_3_ZPOS.txt",net0.n_0_1_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_1_3_ZNEG.txt",net0.n_0_1_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_3_LOCAL.txt",net0.n_0_1_3.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_3_XPOS.txt",net0.n_0_1_3.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_3_XNEG.txt",net0.n_0_1_3.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_3_YPOS.txt",net0.n_0_1_3.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_3_YNEG.txt",net0.n_0_1_3.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_3_ZPOS.txt",net0.n_0_1_3.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_1_3_ZNEG.txt",net0.n_0_1_3.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_0_1_3.txt",net0.n_0_1_3.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_0_LOCAL.txt",net0.n_0_2_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_0_LOCAL.txt",net0.n_0_2_0.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_0_XPOS.txt",net0.n_0_2_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_0_XNEG.txt",net0.n_0_2_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_0_YPOS.txt",net0.n_0_2_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_0_YNEG.txt",net0.n_0_2_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_0_ZPOS.txt",net0.n_0_2_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_0_ZNEG.txt",net0.n_0_2_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_0_LOCAL.txt",net0.n_0_2_0.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_0_XPOS.txt",net0.n_0_2_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_0_XNEG.txt",net0.n_0_2_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_0_YPOS.txt",net0.n_0_2_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_0_YNEG.txt",net0.n_0_2_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_0_ZPOS.txt",net0.n_0_2_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_0_ZNEG.txt",net0.n_0_2_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_0_LOCAL.txt",net0.n_0_2_0.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_0_XPOS.txt",net0.n_0_2_0.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_0_XNEG.txt",net0.n_0_2_0.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_0_YPOS.txt",net0.n_0_2_0.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_0_YNEG.txt",net0.n_0_2_0.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_0_ZPOS.txt",net0.n_0_2_0.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_0_ZNEG.txt",net0.n_0_2_0.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_0_2_0.txt",net0.n_0_2_0.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_1_LOCAL.txt",net0.n_0_2_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_1_LOCAL.txt",net0.n_0_2_1.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_1_XPOS.txt",net0.n_0_2_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_1_XNEG.txt",net0.n_0_2_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_1_YPOS.txt",net0.n_0_2_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_1_YNEG.txt",net0.n_0_2_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_1_ZPOS.txt",net0.n_0_2_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_1_ZNEG.txt",net0.n_0_2_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_1_LOCAL.txt",net0.n_0_2_1.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_1_XPOS.txt",net0.n_0_2_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_1_XNEG.txt",net0.n_0_2_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_1_YPOS.txt",net0.n_0_2_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_1_YNEG.txt",net0.n_0_2_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_1_ZPOS.txt",net0.n_0_2_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_1_ZNEG.txt",net0.n_0_2_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_1_LOCAL.txt",net0.n_0_2_1.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_1_XPOS.txt",net0.n_0_2_1.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_1_XNEG.txt",net0.n_0_2_1.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_1_YPOS.txt",net0.n_0_2_1.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_1_YNEG.txt",net0.n_0_2_1.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_1_ZPOS.txt",net0.n_0_2_1.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_1_ZNEG.txt",net0.n_0_2_1.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_0_2_1.txt",net0.n_0_2_1.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_2_LOCAL.txt",net0.n_0_2_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_2_LOCAL.txt",net0.n_0_2_2.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_2_XPOS.txt",net0.n_0_2_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_2_XNEG.txt",net0.n_0_2_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_2_YPOS.txt",net0.n_0_2_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_2_YNEG.txt",net0.n_0_2_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_2_ZPOS.txt",net0.n_0_2_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_2_ZNEG.txt",net0.n_0_2_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_2_LOCAL.txt",net0.n_0_2_2.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_2_XPOS.txt",net0.n_0_2_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_2_XNEG.txt",net0.n_0_2_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_2_YPOS.txt",net0.n_0_2_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_2_YNEG.txt",net0.n_0_2_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_2_ZPOS.txt",net0.n_0_2_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_2_ZNEG.txt",net0.n_0_2_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_2_LOCAL.txt",net0.n_0_2_2.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_2_XPOS.txt",net0.n_0_2_2.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_2_XNEG.txt",net0.n_0_2_2.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_2_YPOS.txt",net0.n_0_2_2.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_2_YNEG.txt",net0.n_0_2_2.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_2_ZPOS.txt",net0.n_0_2_2.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_2_ZNEG.txt",net0.n_0_2_2.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_0_2_2.txt",net0.n_0_2_2.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_3_LOCAL.txt",net0.n_0_2_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_3_LOCAL.txt",net0.n_0_2_3.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_3_XPOS.txt",net0.n_0_2_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_3_XNEG.txt",net0.n_0_2_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_3_YPOS.txt",net0.n_0_2_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_3_YNEG.txt",net0.n_0_2_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_3_ZPOS.txt",net0.n_0_2_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_2_3_ZNEG.txt",net0.n_0_2_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_3_LOCAL.txt",net0.n_0_2_3.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_3_XPOS.txt",net0.n_0_2_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_3_XNEG.txt",net0.n_0_2_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_3_YPOS.txt",net0.n_0_2_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_3_YNEG.txt",net0.n_0_2_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_3_ZPOS.txt",net0.n_0_2_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_2_3_ZNEG.txt",net0.n_0_2_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_3_LOCAL.txt",net0.n_0_2_3.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_3_XPOS.txt",net0.n_0_2_3.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_3_XNEG.txt",net0.n_0_2_3.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_3_YPOS.txt",net0.n_0_2_3.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_3_YNEG.txt",net0.n_0_2_3.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_3_ZPOS.txt",net0.n_0_2_3.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_2_3_ZNEG.txt",net0.n_0_2_3.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_0_2_3.txt",net0.n_0_2_3.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_0_LOCAL.txt",net0.n_0_3_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_0_LOCAL.txt",net0.n_0_3_0.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_0_XPOS.txt",net0.n_0_3_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_0_XNEG.txt",net0.n_0_3_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_0_YPOS.txt",net0.n_0_3_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_0_YNEG.txt",net0.n_0_3_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_0_ZPOS.txt",net0.n_0_3_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_0_ZNEG.txt",net0.n_0_3_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_0_LOCAL.txt",net0.n_0_3_0.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_0_XPOS.txt",net0.n_0_3_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_0_XNEG.txt",net0.n_0_3_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_0_YPOS.txt",net0.n_0_3_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_0_YNEG.txt",net0.n_0_3_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_0_ZPOS.txt",net0.n_0_3_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_0_ZNEG.txt",net0.n_0_3_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_0_LOCAL.txt",net0.n_0_3_0.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_0_XPOS.txt",net0.n_0_3_0.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_0_XNEG.txt",net0.n_0_3_0.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_0_YPOS.txt",net0.n_0_3_0.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_0_YNEG.txt",net0.n_0_3_0.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_0_ZPOS.txt",net0.n_0_3_0.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_0_ZNEG.txt",net0.n_0_3_0.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_0_3_0.txt",net0.n_0_3_0.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_1_LOCAL.txt",net0.n_0_3_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_1_LOCAL.txt",net0.n_0_3_1.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_1_XPOS.txt",net0.n_0_3_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_1_XNEG.txt",net0.n_0_3_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_1_YPOS.txt",net0.n_0_3_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_1_YNEG.txt",net0.n_0_3_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_1_ZPOS.txt",net0.n_0_3_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_1_ZNEG.txt",net0.n_0_3_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_1_LOCAL.txt",net0.n_0_3_1.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_1_XPOS.txt",net0.n_0_3_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_1_XNEG.txt",net0.n_0_3_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_1_YPOS.txt",net0.n_0_3_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_1_YNEG.txt",net0.n_0_3_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_1_ZPOS.txt",net0.n_0_3_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_1_ZNEG.txt",net0.n_0_3_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_1_LOCAL.txt",net0.n_0_3_1.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_1_XPOS.txt",net0.n_0_3_1.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_1_XNEG.txt",net0.n_0_3_1.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_1_YPOS.txt",net0.n_0_3_1.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_1_YNEG.txt",net0.n_0_3_1.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_1_ZPOS.txt",net0.n_0_3_1.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_1_ZNEG.txt",net0.n_0_3_1.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_0_3_1.txt",net0.n_0_3_1.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_2_LOCAL.txt",net0.n_0_3_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_2_LOCAL.txt",net0.n_0_3_2.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_2_XPOS.txt",net0.n_0_3_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_2_XNEG.txt",net0.n_0_3_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_2_YPOS.txt",net0.n_0_3_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_2_YNEG.txt",net0.n_0_3_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_2_ZPOS.txt",net0.n_0_3_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_2_ZNEG.txt",net0.n_0_3_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_2_LOCAL.txt",net0.n_0_3_2.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_2_XPOS.txt",net0.n_0_3_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_2_XNEG.txt",net0.n_0_3_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_2_YPOS.txt",net0.n_0_3_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_2_YNEG.txt",net0.n_0_3_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_2_ZPOS.txt",net0.n_0_3_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_2_ZNEG.txt",net0.n_0_3_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_2_LOCAL.txt",net0.n_0_3_2.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_2_XPOS.txt",net0.n_0_3_2.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_2_XNEG.txt",net0.n_0_3_2.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_2_YPOS.txt",net0.n_0_3_2.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_2_YNEG.txt",net0.n_0_3_2.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_2_ZPOS.txt",net0.n_0_3_2.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_2_ZNEG.txt",net0.n_0_3_2.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_0_3_2.txt",net0.n_0_3_2.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_3_LOCAL.txt",net0.n_0_3_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_3_LOCAL.txt",net0.n_0_3_3.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_3_XPOS.txt",net0.n_0_3_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_3_XNEG.txt",net0.n_0_3_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_3_YPOS.txt",net0.n_0_3_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_3_YNEG.txt",net0.n_0_3_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_3_ZPOS.txt",net0.n_0_3_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_0_3_3_ZNEG.txt",net0.n_0_3_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_3_LOCAL.txt",net0.n_0_3_3.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_3_XPOS.txt",net0.n_0_3_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_3_XNEG.txt",net0.n_0_3_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_3_YPOS.txt",net0.n_0_3_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_3_YNEG.txt",net0.n_0_3_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_3_ZPOS.txt",net0.n_0_3_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_0_3_3_ZNEG.txt",net0.n_0_3_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_3_LOCAL.txt",net0.n_0_3_3.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_3_XPOS.txt",net0.n_0_3_3.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_3_XNEG.txt",net0.n_0_3_3.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_3_YPOS.txt",net0.n_0_3_3.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_3_YNEG.txt",net0.n_0_3_3.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_3_ZPOS.txt",net0.n_0_3_3.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_0_3_3_ZNEG.txt",net0.n_0_3_3.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_0_3_3.txt",net0.n_0_3_3.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_0_LOCAL.txt",net0.n_1_0_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_0_LOCAL.txt",net0.n_1_0_0.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_0_XPOS.txt",net0.n_1_0_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_0_XNEG.txt",net0.n_1_0_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_0_YPOS.txt",net0.n_1_0_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_0_YNEG.txt",net0.n_1_0_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_0_ZPOS.txt",net0.n_1_0_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_0_ZNEG.txt",net0.n_1_0_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_0_LOCAL.txt",net0.n_1_0_0.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_0_XPOS.txt",net0.n_1_0_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_0_XNEG.txt",net0.n_1_0_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_0_YPOS.txt",net0.n_1_0_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_0_YNEG.txt",net0.n_1_0_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_0_ZPOS.txt",net0.n_1_0_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_0_ZNEG.txt",net0.n_1_0_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_0_LOCAL.txt",net0.n_1_0_0.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_0_XPOS.txt",net0.n_1_0_0.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_0_XNEG.txt",net0.n_1_0_0.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_0_YPOS.txt",net0.n_1_0_0.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_0_YNEG.txt",net0.n_1_0_0.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_0_ZPOS.txt",net0.n_1_0_0.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_0_ZNEG.txt",net0.n_1_0_0.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_1_0_0.txt",net0.n_1_0_0.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_1_LOCAL.txt",net0.n_1_0_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_1_LOCAL.txt",net0.n_1_0_1.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_1_XPOS.txt",net0.n_1_0_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_1_XNEG.txt",net0.n_1_0_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_1_YPOS.txt",net0.n_1_0_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_1_YNEG.txt",net0.n_1_0_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_1_ZPOS.txt",net0.n_1_0_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_1_ZNEG.txt",net0.n_1_0_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_1_LOCAL.txt",net0.n_1_0_1.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_1_XPOS.txt",net0.n_1_0_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_1_XNEG.txt",net0.n_1_0_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_1_YPOS.txt",net0.n_1_0_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_1_YNEG.txt",net0.n_1_0_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_1_ZPOS.txt",net0.n_1_0_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_1_ZNEG.txt",net0.n_1_0_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_1_LOCAL.txt",net0.n_1_0_1.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_1_XPOS.txt",net0.n_1_0_1.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_1_XNEG.txt",net0.n_1_0_1.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_1_YPOS.txt",net0.n_1_0_1.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_1_YNEG.txt",net0.n_1_0_1.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_1_ZPOS.txt",net0.n_1_0_1.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_1_ZNEG.txt",net0.n_1_0_1.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_1_0_1.txt",net0.n_1_0_1.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_2_LOCAL.txt",net0.n_1_0_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_2_LOCAL.txt",net0.n_1_0_2.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_2_XPOS.txt",net0.n_1_0_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_2_XNEG.txt",net0.n_1_0_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_2_YPOS.txt",net0.n_1_0_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_2_YNEG.txt",net0.n_1_0_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_2_ZPOS.txt",net0.n_1_0_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_2_ZNEG.txt",net0.n_1_0_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_2_LOCAL.txt",net0.n_1_0_2.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_2_XPOS.txt",net0.n_1_0_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_2_XNEG.txt",net0.n_1_0_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_2_YPOS.txt",net0.n_1_0_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_2_YNEG.txt",net0.n_1_0_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_2_ZPOS.txt",net0.n_1_0_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_2_ZNEG.txt",net0.n_1_0_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_2_LOCAL.txt",net0.n_1_0_2.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_2_XPOS.txt",net0.n_1_0_2.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_2_XNEG.txt",net0.n_1_0_2.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_2_YPOS.txt",net0.n_1_0_2.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_2_YNEG.txt",net0.n_1_0_2.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_2_ZPOS.txt",net0.n_1_0_2.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_2_ZNEG.txt",net0.n_1_0_2.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_1_0_2.txt",net0.n_1_0_2.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_3_LOCAL.txt",net0.n_1_0_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_3_LOCAL.txt",net0.n_1_0_3.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_3_XPOS.txt",net0.n_1_0_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_3_XNEG.txt",net0.n_1_0_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_3_YPOS.txt",net0.n_1_0_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_3_YNEG.txt",net0.n_1_0_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_3_ZPOS.txt",net0.n_1_0_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_0_3_ZNEG.txt",net0.n_1_0_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_3_LOCAL.txt",net0.n_1_0_3.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_3_XPOS.txt",net0.n_1_0_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_3_XNEG.txt",net0.n_1_0_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_3_YPOS.txt",net0.n_1_0_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_3_YNEG.txt",net0.n_1_0_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_3_ZPOS.txt",net0.n_1_0_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_0_3_ZNEG.txt",net0.n_1_0_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_3_LOCAL.txt",net0.n_1_0_3.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_3_XPOS.txt",net0.n_1_0_3.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_3_XNEG.txt",net0.n_1_0_3.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_3_YPOS.txt",net0.n_1_0_3.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_3_YNEG.txt",net0.n_1_0_3.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_3_ZPOS.txt",net0.n_1_0_3.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_0_3_ZNEG.txt",net0.n_1_0_3.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_1_0_3.txt",net0.n_1_0_3.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_0_LOCAL.txt",net0.n_1_1_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_0_LOCAL.txt",net0.n_1_1_0.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_0_XPOS.txt",net0.n_1_1_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_0_XNEG.txt",net0.n_1_1_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_0_YPOS.txt",net0.n_1_1_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_0_YNEG.txt",net0.n_1_1_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_0_ZPOS.txt",net0.n_1_1_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_0_ZNEG.txt",net0.n_1_1_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_0_LOCAL.txt",net0.n_1_1_0.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_0_XPOS.txt",net0.n_1_1_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_0_XNEG.txt",net0.n_1_1_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_0_YPOS.txt",net0.n_1_1_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_0_YNEG.txt",net0.n_1_1_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_0_ZPOS.txt",net0.n_1_1_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_0_ZNEG.txt",net0.n_1_1_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_0_LOCAL.txt",net0.n_1_1_0.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_0_XPOS.txt",net0.n_1_1_0.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_0_XNEG.txt",net0.n_1_1_0.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_0_YPOS.txt",net0.n_1_1_0.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_0_YNEG.txt",net0.n_1_1_0.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_0_ZPOS.txt",net0.n_1_1_0.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_0_ZNEG.txt",net0.n_1_1_0.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_1_1_0.txt",net0.n_1_1_0.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_1_LOCAL.txt",net0.n_1_1_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_1_LOCAL.txt",net0.n_1_1_1.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_1_XPOS.txt",net0.n_1_1_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_1_XNEG.txt",net0.n_1_1_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_1_YPOS.txt",net0.n_1_1_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_1_YNEG.txt",net0.n_1_1_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_1_ZPOS.txt",net0.n_1_1_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_1_ZNEG.txt",net0.n_1_1_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_1_LOCAL.txt",net0.n_1_1_1.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_1_XPOS.txt",net0.n_1_1_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_1_XNEG.txt",net0.n_1_1_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_1_YPOS.txt",net0.n_1_1_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_1_YNEG.txt",net0.n_1_1_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_1_ZPOS.txt",net0.n_1_1_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_1_ZNEG.txt",net0.n_1_1_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_1_LOCAL.txt",net0.n_1_1_1.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_1_XPOS.txt",net0.n_1_1_1.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_1_XNEG.txt",net0.n_1_1_1.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_1_YPOS.txt",net0.n_1_1_1.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_1_YNEG.txt",net0.n_1_1_1.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_1_ZPOS.txt",net0.n_1_1_1.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_1_ZNEG.txt",net0.n_1_1_1.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_1_1_1.txt",net0.n_1_1_1.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_2_LOCAL.txt",net0.n_1_1_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_2_LOCAL.txt",net0.n_1_1_2.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_2_XPOS.txt",net0.n_1_1_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_2_XNEG.txt",net0.n_1_1_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_2_YPOS.txt",net0.n_1_1_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_2_YNEG.txt",net0.n_1_1_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_2_ZPOS.txt",net0.n_1_1_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_2_ZNEG.txt",net0.n_1_1_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_2_LOCAL.txt",net0.n_1_1_2.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_2_XPOS.txt",net0.n_1_1_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_2_XNEG.txt",net0.n_1_1_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_2_YPOS.txt",net0.n_1_1_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_2_YNEG.txt",net0.n_1_1_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_2_ZPOS.txt",net0.n_1_1_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_2_ZNEG.txt",net0.n_1_1_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_2_LOCAL.txt",net0.n_1_1_2.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_2_XPOS.txt",net0.n_1_1_2.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_2_XNEG.txt",net0.n_1_1_2.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_2_YPOS.txt",net0.n_1_1_2.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_2_YNEG.txt",net0.n_1_1_2.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_2_ZPOS.txt",net0.n_1_1_2.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_2_ZNEG.txt",net0.n_1_1_2.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_1_1_2.txt",net0.n_1_1_2.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_3_LOCAL.txt",net0.n_1_1_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_3_LOCAL.txt",net0.n_1_1_3.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_3_XPOS.txt",net0.n_1_1_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_3_XNEG.txt",net0.n_1_1_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_3_YPOS.txt",net0.n_1_1_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_3_YNEG.txt",net0.n_1_1_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_3_ZPOS.txt",net0.n_1_1_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_1_3_ZNEG.txt",net0.n_1_1_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_3_LOCAL.txt",net0.n_1_1_3.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_3_XPOS.txt",net0.n_1_1_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_3_XNEG.txt",net0.n_1_1_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_3_YPOS.txt",net0.n_1_1_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_3_YNEG.txt",net0.n_1_1_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_3_ZPOS.txt",net0.n_1_1_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_1_3_ZNEG.txt",net0.n_1_1_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_3_LOCAL.txt",net0.n_1_1_3.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_3_XPOS.txt",net0.n_1_1_3.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_3_XNEG.txt",net0.n_1_1_3.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_3_YPOS.txt",net0.n_1_1_3.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_3_YNEG.txt",net0.n_1_1_3.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_3_ZPOS.txt",net0.n_1_1_3.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_1_3_ZNEG.txt",net0.n_1_1_3.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_1_1_3.txt",net0.n_1_1_3.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_0_LOCAL.txt",net0.n_1_2_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_0_LOCAL.txt",net0.n_1_2_0.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_0_XPOS.txt",net0.n_1_2_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_0_XNEG.txt",net0.n_1_2_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_0_YPOS.txt",net0.n_1_2_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_0_YNEG.txt",net0.n_1_2_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_0_ZPOS.txt",net0.n_1_2_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_0_ZNEG.txt",net0.n_1_2_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_0_LOCAL.txt",net0.n_1_2_0.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_0_XPOS.txt",net0.n_1_2_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_0_XNEG.txt",net0.n_1_2_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_0_YPOS.txt",net0.n_1_2_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_0_YNEG.txt",net0.n_1_2_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_0_ZPOS.txt",net0.n_1_2_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_0_ZNEG.txt",net0.n_1_2_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_0_LOCAL.txt",net0.n_1_2_0.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_0_XPOS.txt",net0.n_1_2_0.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_0_XNEG.txt",net0.n_1_2_0.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_0_YPOS.txt",net0.n_1_2_0.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_0_YNEG.txt",net0.n_1_2_0.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_0_ZPOS.txt",net0.n_1_2_0.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_0_ZNEG.txt",net0.n_1_2_0.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_1_2_0.txt",net0.n_1_2_0.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_1_LOCAL.txt",net0.n_1_2_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_1_LOCAL.txt",net0.n_1_2_1.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_1_XPOS.txt",net0.n_1_2_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_1_XNEG.txt",net0.n_1_2_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_1_YPOS.txt",net0.n_1_2_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_1_YNEG.txt",net0.n_1_2_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_1_ZPOS.txt",net0.n_1_2_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_1_ZNEG.txt",net0.n_1_2_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_1_LOCAL.txt",net0.n_1_2_1.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_1_XPOS.txt",net0.n_1_2_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_1_XNEG.txt",net0.n_1_2_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_1_YPOS.txt",net0.n_1_2_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_1_YNEG.txt",net0.n_1_2_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_1_ZPOS.txt",net0.n_1_2_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_1_ZNEG.txt",net0.n_1_2_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_1_LOCAL.txt",net0.n_1_2_1.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_1_XPOS.txt",net0.n_1_2_1.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_1_XNEG.txt",net0.n_1_2_1.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_1_YPOS.txt",net0.n_1_2_1.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_1_YNEG.txt",net0.n_1_2_1.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_1_ZPOS.txt",net0.n_1_2_1.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_1_ZNEG.txt",net0.n_1_2_1.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_1_2_1.txt",net0.n_1_2_1.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_2_LOCAL.txt",net0.n_1_2_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_2_LOCAL.txt",net0.n_1_2_2.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_2_XPOS.txt",net0.n_1_2_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_2_XNEG.txt",net0.n_1_2_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_2_YPOS.txt",net0.n_1_2_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_2_YNEG.txt",net0.n_1_2_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_2_ZPOS.txt",net0.n_1_2_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_2_ZNEG.txt",net0.n_1_2_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_2_LOCAL.txt",net0.n_1_2_2.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_2_XPOS.txt",net0.n_1_2_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_2_XNEG.txt",net0.n_1_2_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_2_YPOS.txt",net0.n_1_2_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_2_YNEG.txt",net0.n_1_2_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_2_ZPOS.txt",net0.n_1_2_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_2_ZNEG.txt",net0.n_1_2_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_2_LOCAL.txt",net0.n_1_2_2.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_2_XPOS.txt",net0.n_1_2_2.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_2_XNEG.txt",net0.n_1_2_2.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_2_YPOS.txt",net0.n_1_2_2.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_2_YNEG.txt",net0.n_1_2_2.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_2_ZPOS.txt",net0.n_1_2_2.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_2_ZNEG.txt",net0.n_1_2_2.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_1_2_2.txt",net0.n_1_2_2.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_3_LOCAL.txt",net0.n_1_2_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_3_LOCAL.txt",net0.n_1_2_3.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_3_XPOS.txt",net0.n_1_2_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_3_XNEG.txt",net0.n_1_2_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_3_YPOS.txt",net0.n_1_2_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_3_YNEG.txt",net0.n_1_2_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_3_ZPOS.txt",net0.n_1_2_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_2_3_ZNEG.txt",net0.n_1_2_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_3_LOCAL.txt",net0.n_1_2_3.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_3_XPOS.txt",net0.n_1_2_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_3_XNEG.txt",net0.n_1_2_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_3_YPOS.txt",net0.n_1_2_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_3_YNEG.txt",net0.n_1_2_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_3_ZPOS.txt",net0.n_1_2_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_2_3_ZNEG.txt",net0.n_1_2_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_3_LOCAL.txt",net0.n_1_2_3.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_3_XPOS.txt",net0.n_1_2_3.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_3_XNEG.txt",net0.n_1_2_3.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_3_YPOS.txt",net0.n_1_2_3.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_3_YNEG.txt",net0.n_1_2_3.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_3_ZPOS.txt",net0.n_1_2_3.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_2_3_ZNEG.txt",net0.n_1_2_3.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_1_2_3.txt",net0.n_1_2_3.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_0_LOCAL.txt",net0.n_1_3_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_0_LOCAL.txt",net0.n_1_3_0.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_0_XPOS.txt",net0.n_1_3_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_0_XNEG.txt",net0.n_1_3_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_0_YPOS.txt",net0.n_1_3_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_0_YNEG.txt",net0.n_1_3_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_0_ZPOS.txt",net0.n_1_3_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_0_ZNEG.txt",net0.n_1_3_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_0_LOCAL.txt",net0.n_1_3_0.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_0_XPOS.txt",net0.n_1_3_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_0_XNEG.txt",net0.n_1_3_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_0_YPOS.txt",net0.n_1_3_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_0_YNEG.txt",net0.n_1_3_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_0_ZPOS.txt",net0.n_1_3_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_0_ZNEG.txt",net0.n_1_3_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_0_LOCAL.txt",net0.n_1_3_0.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_0_XPOS.txt",net0.n_1_3_0.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_0_XNEG.txt",net0.n_1_3_0.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_0_YPOS.txt",net0.n_1_3_0.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_0_YNEG.txt",net0.n_1_3_0.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_0_ZPOS.txt",net0.n_1_3_0.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_0_ZNEG.txt",net0.n_1_3_0.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_1_3_0.txt",net0.n_1_3_0.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_1_LOCAL.txt",net0.n_1_3_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_1_LOCAL.txt",net0.n_1_3_1.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_1_XPOS.txt",net0.n_1_3_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_1_XNEG.txt",net0.n_1_3_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_1_YPOS.txt",net0.n_1_3_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_1_YNEG.txt",net0.n_1_3_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_1_ZPOS.txt",net0.n_1_3_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_1_ZNEG.txt",net0.n_1_3_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_1_LOCAL.txt",net0.n_1_3_1.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_1_XPOS.txt",net0.n_1_3_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_1_XNEG.txt",net0.n_1_3_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_1_YPOS.txt",net0.n_1_3_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_1_YNEG.txt",net0.n_1_3_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_1_ZPOS.txt",net0.n_1_3_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_1_ZNEG.txt",net0.n_1_3_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_1_LOCAL.txt",net0.n_1_3_1.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_1_XPOS.txt",net0.n_1_3_1.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_1_XNEG.txt",net0.n_1_3_1.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_1_YPOS.txt",net0.n_1_3_1.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_1_YNEG.txt",net0.n_1_3_1.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_1_ZPOS.txt",net0.n_1_3_1.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_1_ZNEG.txt",net0.n_1_3_1.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_1_3_1.txt",net0.n_1_3_1.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_2_LOCAL.txt",net0.n_1_3_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_2_LOCAL.txt",net0.n_1_3_2.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_2_XPOS.txt",net0.n_1_3_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_2_XNEG.txt",net0.n_1_3_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_2_YPOS.txt",net0.n_1_3_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_2_YNEG.txt",net0.n_1_3_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_2_ZPOS.txt",net0.n_1_3_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_2_ZNEG.txt",net0.n_1_3_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_2_LOCAL.txt",net0.n_1_3_2.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_2_XPOS.txt",net0.n_1_3_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_2_XNEG.txt",net0.n_1_3_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_2_YPOS.txt",net0.n_1_3_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_2_YNEG.txt",net0.n_1_3_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_2_ZPOS.txt",net0.n_1_3_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_2_ZNEG.txt",net0.n_1_3_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_2_LOCAL.txt",net0.n_1_3_2.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_2_XPOS.txt",net0.n_1_3_2.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_2_XNEG.txt",net0.n_1_3_2.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_2_YPOS.txt",net0.n_1_3_2.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_2_YNEG.txt",net0.n_1_3_2.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_2_ZPOS.txt",net0.n_1_3_2.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_2_ZNEG.txt",net0.n_1_3_2.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_1_3_2.txt",net0.n_1_3_2.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_3_LOCAL.txt",net0.n_1_3_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_3_LOCAL.txt",net0.n_1_3_3.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_3_XPOS.txt",net0.n_1_3_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_3_XNEG.txt",net0.n_1_3_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_3_YPOS.txt",net0.n_1_3_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_3_YNEG.txt",net0.n_1_3_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_3_ZPOS.txt",net0.n_1_3_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_1_3_3_ZNEG.txt",net0.n_1_3_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_3_LOCAL.txt",net0.n_1_3_3.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_3_XPOS.txt",net0.n_1_3_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_3_XNEG.txt",net0.n_1_3_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_3_YPOS.txt",net0.n_1_3_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_3_YNEG.txt",net0.n_1_3_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_3_ZPOS.txt",net0.n_1_3_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_1_3_3_ZNEG.txt",net0.n_1_3_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_3_LOCAL.txt",net0.n_1_3_3.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_3_XPOS.txt",net0.n_1_3_3.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_3_XNEG.txt",net0.n_1_3_3.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_3_YPOS.txt",net0.n_1_3_3.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_3_YNEG.txt",net0.n_1_3_3.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_3_ZPOS.txt",net0.n_1_3_3.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_1_3_3_ZNEG.txt",net0.n_1_3_3.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_1_3_3.txt",net0.n_1_3_3.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_0_LOCAL.txt",net0.n_2_0_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_0_LOCAL.txt",net0.n_2_0_0.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_0_XPOS.txt",net0.n_2_0_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_0_XNEG.txt",net0.n_2_0_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_0_YPOS.txt",net0.n_2_0_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_0_YNEG.txt",net0.n_2_0_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_0_ZPOS.txt",net0.n_2_0_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_0_ZNEG.txt",net0.n_2_0_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_0_LOCAL.txt",net0.n_2_0_0.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_0_XPOS.txt",net0.n_2_0_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_0_XNEG.txt",net0.n_2_0_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_0_YPOS.txt",net0.n_2_0_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_0_YNEG.txt",net0.n_2_0_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_0_ZPOS.txt",net0.n_2_0_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_0_ZNEG.txt",net0.n_2_0_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_0_LOCAL.txt",net0.n_2_0_0.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_0_XPOS.txt",net0.n_2_0_0.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_0_XNEG.txt",net0.n_2_0_0.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_0_YPOS.txt",net0.n_2_0_0.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_0_YNEG.txt",net0.n_2_0_0.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_0_ZPOS.txt",net0.n_2_0_0.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_0_ZNEG.txt",net0.n_2_0_0.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_2_0_0.txt",net0.n_2_0_0.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_1_LOCAL.txt",net0.n_2_0_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_1_LOCAL.txt",net0.n_2_0_1.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_1_XPOS.txt",net0.n_2_0_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_1_XNEG.txt",net0.n_2_0_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_1_YPOS.txt",net0.n_2_0_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_1_YNEG.txt",net0.n_2_0_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_1_ZPOS.txt",net0.n_2_0_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_1_ZNEG.txt",net0.n_2_0_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_1_LOCAL.txt",net0.n_2_0_1.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_1_XPOS.txt",net0.n_2_0_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_1_XNEG.txt",net0.n_2_0_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_1_YPOS.txt",net0.n_2_0_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_1_YNEG.txt",net0.n_2_0_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_1_ZPOS.txt",net0.n_2_0_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_1_ZNEG.txt",net0.n_2_0_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_1_LOCAL.txt",net0.n_2_0_1.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_1_XPOS.txt",net0.n_2_0_1.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_1_XNEG.txt",net0.n_2_0_1.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_1_YPOS.txt",net0.n_2_0_1.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_1_YNEG.txt",net0.n_2_0_1.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_1_ZPOS.txt",net0.n_2_0_1.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_1_ZNEG.txt",net0.n_2_0_1.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_2_0_1.txt",net0.n_2_0_1.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_2_LOCAL.txt",net0.n_2_0_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_2_LOCAL.txt",net0.n_2_0_2.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_2_XPOS.txt",net0.n_2_0_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_2_XNEG.txt",net0.n_2_0_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_2_YPOS.txt",net0.n_2_0_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_2_YNEG.txt",net0.n_2_0_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_2_ZPOS.txt",net0.n_2_0_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_2_ZNEG.txt",net0.n_2_0_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_2_LOCAL.txt",net0.n_2_0_2.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_2_XPOS.txt",net0.n_2_0_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_2_XNEG.txt",net0.n_2_0_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_2_YPOS.txt",net0.n_2_0_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_2_YNEG.txt",net0.n_2_0_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_2_ZPOS.txt",net0.n_2_0_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_2_ZNEG.txt",net0.n_2_0_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_2_LOCAL.txt",net0.n_2_0_2.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_2_XPOS.txt",net0.n_2_0_2.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_2_XNEG.txt",net0.n_2_0_2.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_2_YPOS.txt",net0.n_2_0_2.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_2_YNEG.txt",net0.n_2_0_2.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_2_ZPOS.txt",net0.n_2_0_2.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_2_ZNEG.txt",net0.n_2_0_2.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_2_0_2.txt",net0.n_2_0_2.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_3_LOCAL.txt",net0.n_2_0_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_3_LOCAL.txt",net0.n_2_0_3.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_3_XPOS.txt",net0.n_2_0_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_3_XNEG.txt",net0.n_2_0_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_3_YPOS.txt",net0.n_2_0_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_3_YNEG.txt",net0.n_2_0_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_3_ZPOS.txt",net0.n_2_0_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_0_3_ZNEG.txt",net0.n_2_0_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_3_LOCAL.txt",net0.n_2_0_3.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_3_XPOS.txt",net0.n_2_0_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_3_XNEG.txt",net0.n_2_0_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_3_YPOS.txt",net0.n_2_0_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_3_YNEG.txt",net0.n_2_0_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_3_ZPOS.txt",net0.n_2_0_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_0_3_ZNEG.txt",net0.n_2_0_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_3_LOCAL.txt",net0.n_2_0_3.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_3_XPOS.txt",net0.n_2_0_3.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_3_XNEG.txt",net0.n_2_0_3.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_3_YPOS.txt",net0.n_2_0_3.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_3_YNEG.txt",net0.n_2_0_3.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_3_ZPOS.txt",net0.n_2_0_3.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_0_3_ZNEG.txt",net0.n_2_0_3.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_2_0_3.txt",net0.n_2_0_3.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_0_LOCAL.txt",net0.n_2_1_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_0_LOCAL.txt",net0.n_2_1_0.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_0_XPOS.txt",net0.n_2_1_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_0_XNEG.txt",net0.n_2_1_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_0_YPOS.txt",net0.n_2_1_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_0_YNEG.txt",net0.n_2_1_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_0_ZPOS.txt",net0.n_2_1_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_0_ZNEG.txt",net0.n_2_1_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_0_LOCAL.txt",net0.n_2_1_0.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_0_XPOS.txt",net0.n_2_1_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_0_XNEG.txt",net0.n_2_1_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_0_YPOS.txt",net0.n_2_1_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_0_YNEG.txt",net0.n_2_1_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_0_ZPOS.txt",net0.n_2_1_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_0_ZNEG.txt",net0.n_2_1_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_0_LOCAL.txt",net0.n_2_1_0.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_0_XPOS.txt",net0.n_2_1_0.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_0_XNEG.txt",net0.n_2_1_0.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_0_YPOS.txt",net0.n_2_1_0.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_0_YNEG.txt",net0.n_2_1_0.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_0_ZPOS.txt",net0.n_2_1_0.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_0_ZNEG.txt",net0.n_2_1_0.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_2_1_0.txt",net0.n_2_1_0.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_1_LOCAL.txt",net0.n_2_1_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_1_LOCAL.txt",net0.n_2_1_1.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_1_XPOS.txt",net0.n_2_1_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_1_XNEG.txt",net0.n_2_1_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_1_YPOS.txt",net0.n_2_1_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_1_YNEG.txt",net0.n_2_1_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_1_ZPOS.txt",net0.n_2_1_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_1_ZNEG.txt",net0.n_2_1_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_1_LOCAL.txt",net0.n_2_1_1.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_1_XPOS.txt",net0.n_2_1_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_1_XNEG.txt",net0.n_2_1_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_1_YPOS.txt",net0.n_2_1_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_1_YNEG.txt",net0.n_2_1_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_1_ZPOS.txt",net0.n_2_1_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_1_ZNEG.txt",net0.n_2_1_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_1_LOCAL.txt",net0.n_2_1_1.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_1_XPOS.txt",net0.n_2_1_1.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_1_XNEG.txt",net0.n_2_1_1.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_1_YPOS.txt",net0.n_2_1_1.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_1_YNEG.txt",net0.n_2_1_1.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_1_ZPOS.txt",net0.n_2_1_1.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_1_ZNEG.txt",net0.n_2_1_1.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_2_1_1.txt",net0.n_2_1_1.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_2_LOCAL.txt",net0.n_2_1_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_2_LOCAL.txt",net0.n_2_1_2.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_2_XPOS.txt",net0.n_2_1_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_2_XNEG.txt",net0.n_2_1_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_2_YPOS.txt",net0.n_2_1_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_2_YNEG.txt",net0.n_2_1_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_2_ZPOS.txt",net0.n_2_1_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_2_ZNEG.txt",net0.n_2_1_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_2_LOCAL.txt",net0.n_2_1_2.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_2_XPOS.txt",net0.n_2_1_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_2_XNEG.txt",net0.n_2_1_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_2_YPOS.txt",net0.n_2_1_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_2_YNEG.txt",net0.n_2_1_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_2_ZPOS.txt",net0.n_2_1_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_2_ZNEG.txt",net0.n_2_1_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_2_LOCAL.txt",net0.n_2_1_2.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_2_XPOS.txt",net0.n_2_1_2.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_2_XNEG.txt",net0.n_2_1_2.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_2_YPOS.txt",net0.n_2_1_2.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_2_YNEG.txt",net0.n_2_1_2.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_2_ZPOS.txt",net0.n_2_1_2.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_2_ZNEG.txt",net0.n_2_1_2.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_2_1_2.txt",net0.n_2_1_2.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_3_LOCAL.txt",net0.n_2_1_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_3_LOCAL.txt",net0.n_2_1_3.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_3_XPOS.txt",net0.n_2_1_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_3_XNEG.txt",net0.n_2_1_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_3_YPOS.txt",net0.n_2_1_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_3_YNEG.txt",net0.n_2_1_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_3_ZPOS.txt",net0.n_2_1_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_1_3_ZNEG.txt",net0.n_2_1_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_3_LOCAL.txt",net0.n_2_1_3.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_3_XPOS.txt",net0.n_2_1_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_3_XNEG.txt",net0.n_2_1_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_3_YPOS.txt",net0.n_2_1_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_3_YNEG.txt",net0.n_2_1_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_3_ZPOS.txt",net0.n_2_1_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_1_3_ZNEG.txt",net0.n_2_1_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_3_LOCAL.txt",net0.n_2_1_3.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_3_XPOS.txt",net0.n_2_1_3.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_3_XNEG.txt",net0.n_2_1_3.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_3_YPOS.txt",net0.n_2_1_3.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_3_YNEG.txt",net0.n_2_1_3.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_3_ZPOS.txt",net0.n_2_1_3.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_1_3_ZNEG.txt",net0.n_2_1_3.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_2_1_3.txt",net0.n_2_1_3.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_0_LOCAL.txt",net0.n_2_2_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_0_LOCAL.txt",net0.n_2_2_0.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_0_XPOS.txt",net0.n_2_2_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_0_XNEG.txt",net0.n_2_2_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_0_YPOS.txt",net0.n_2_2_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_0_YNEG.txt",net0.n_2_2_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_0_ZPOS.txt",net0.n_2_2_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_0_ZNEG.txt",net0.n_2_2_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_0_LOCAL.txt",net0.n_2_2_0.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_0_XPOS.txt",net0.n_2_2_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_0_XNEG.txt",net0.n_2_2_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_0_YPOS.txt",net0.n_2_2_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_0_YNEG.txt",net0.n_2_2_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_0_ZPOS.txt",net0.n_2_2_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_0_ZNEG.txt",net0.n_2_2_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_0_LOCAL.txt",net0.n_2_2_0.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_0_XPOS.txt",net0.n_2_2_0.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_0_XNEG.txt",net0.n_2_2_0.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_0_YPOS.txt",net0.n_2_2_0.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_0_YNEG.txt",net0.n_2_2_0.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_0_ZPOS.txt",net0.n_2_2_0.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_0_ZNEG.txt",net0.n_2_2_0.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_2_2_0.txt",net0.n_2_2_0.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_1_LOCAL.txt",net0.n_2_2_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_1_LOCAL.txt",net0.n_2_2_1.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_1_XPOS.txt",net0.n_2_2_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_1_XNEG.txt",net0.n_2_2_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_1_YPOS.txt",net0.n_2_2_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_1_YNEG.txt",net0.n_2_2_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_1_ZPOS.txt",net0.n_2_2_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_1_ZNEG.txt",net0.n_2_2_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_1_LOCAL.txt",net0.n_2_2_1.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_1_XPOS.txt",net0.n_2_2_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_1_XNEG.txt",net0.n_2_2_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_1_YPOS.txt",net0.n_2_2_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_1_YNEG.txt",net0.n_2_2_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_1_ZPOS.txt",net0.n_2_2_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_1_ZNEG.txt",net0.n_2_2_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_1_LOCAL.txt",net0.n_2_2_1.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_1_XPOS.txt",net0.n_2_2_1.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_1_XNEG.txt",net0.n_2_2_1.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_1_YPOS.txt",net0.n_2_2_1.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_1_YNEG.txt",net0.n_2_2_1.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_1_ZPOS.txt",net0.n_2_2_1.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_1_ZNEG.txt",net0.n_2_2_1.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_2_2_1.txt",net0.n_2_2_1.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_2_LOCAL.txt",net0.n_2_2_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_2_LOCAL.txt",net0.n_2_2_2.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_2_XPOS.txt",net0.n_2_2_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_2_XNEG.txt",net0.n_2_2_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_2_YPOS.txt",net0.n_2_2_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_2_YNEG.txt",net0.n_2_2_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_2_ZPOS.txt",net0.n_2_2_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_2_ZNEG.txt",net0.n_2_2_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_2_LOCAL.txt",net0.n_2_2_2.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_2_XPOS.txt",net0.n_2_2_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_2_XNEG.txt",net0.n_2_2_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_2_YPOS.txt",net0.n_2_2_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_2_YNEG.txt",net0.n_2_2_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_2_ZPOS.txt",net0.n_2_2_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_2_ZNEG.txt",net0.n_2_2_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_2_LOCAL.txt",net0.n_2_2_2.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_2_XPOS.txt",net0.n_2_2_2.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_2_XNEG.txt",net0.n_2_2_2.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_2_YPOS.txt",net0.n_2_2_2.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_2_YNEG.txt",net0.n_2_2_2.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_2_ZPOS.txt",net0.n_2_2_2.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_2_ZNEG.txt",net0.n_2_2_2.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_2_2_2.txt",net0.n_2_2_2.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_3_LOCAL.txt",net0.n_2_2_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_3_LOCAL.txt",net0.n_2_2_3.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_3_XPOS.txt",net0.n_2_2_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_3_XNEG.txt",net0.n_2_2_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_3_YPOS.txt",net0.n_2_2_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_3_YNEG.txt",net0.n_2_2_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_3_ZPOS.txt",net0.n_2_2_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_2_3_ZNEG.txt",net0.n_2_2_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_3_LOCAL.txt",net0.n_2_2_3.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_3_XPOS.txt",net0.n_2_2_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_3_XNEG.txt",net0.n_2_2_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_3_YPOS.txt",net0.n_2_2_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_3_YNEG.txt",net0.n_2_2_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_3_ZPOS.txt",net0.n_2_2_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_2_3_ZNEG.txt",net0.n_2_2_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_3_LOCAL.txt",net0.n_2_2_3.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_3_XPOS.txt",net0.n_2_2_3.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_3_XNEG.txt",net0.n_2_2_3.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_3_YPOS.txt",net0.n_2_2_3.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_3_YNEG.txt",net0.n_2_2_3.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_3_ZPOS.txt",net0.n_2_2_3.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_2_3_ZNEG.txt",net0.n_2_2_3.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_2_2_3.txt",net0.n_2_2_3.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_0_LOCAL.txt",net0.n_2_3_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_0_LOCAL.txt",net0.n_2_3_0.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_0_XPOS.txt",net0.n_2_3_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_0_XNEG.txt",net0.n_2_3_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_0_YPOS.txt",net0.n_2_3_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_0_YNEG.txt",net0.n_2_3_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_0_ZPOS.txt",net0.n_2_3_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_0_ZNEG.txt",net0.n_2_3_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_0_LOCAL.txt",net0.n_2_3_0.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_0_XPOS.txt",net0.n_2_3_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_0_XNEG.txt",net0.n_2_3_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_0_YPOS.txt",net0.n_2_3_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_0_YNEG.txt",net0.n_2_3_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_0_ZPOS.txt",net0.n_2_3_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_0_ZNEG.txt",net0.n_2_3_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_0_LOCAL.txt",net0.n_2_3_0.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_0_XPOS.txt",net0.n_2_3_0.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_0_XNEG.txt",net0.n_2_3_0.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_0_YPOS.txt",net0.n_2_3_0.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_0_YNEG.txt",net0.n_2_3_0.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_0_ZPOS.txt",net0.n_2_3_0.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_0_ZNEG.txt",net0.n_2_3_0.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_2_3_0.txt",net0.n_2_3_0.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_1_LOCAL.txt",net0.n_2_3_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_1_LOCAL.txt",net0.n_2_3_1.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_1_XPOS.txt",net0.n_2_3_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_1_XNEG.txt",net0.n_2_3_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_1_YPOS.txt",net0.n_2_3_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_1_YNEG.txt",net0.n_2_3_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_1_ZPOS.txt",net0.n_2_3_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_1_ZNEG.txt",net0.n_2_3_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_1_LOCAL.txt",net0.n_2_3_1.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_1_XPOS.txt",net0.n_2_3_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_1_XNEG.txt",net0.n_2_3_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_1_YPOS.txt",net0.n_2_3_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_1_YNEG.txt",net0.n_2_3_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_1_ZPOS.txt",net0.n_2_3_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_1_ZNEG.txt",net0.n_2_3_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_1_LOCAL.txt",net0.n_2_3_1.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_1_XPOS.txt",net0.n_2_3_1.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_1_XNEG.txt",net0.n_2_3_1.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_1_YPOS.txt",net0.n_2_3_1.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_1_YNEG.txt",net0.n_2_3_1.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_1_ZPOS.txt",net0.n_2_3_1.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_1_ZNEG.txt",net0.n_2_3_1.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_2_3_1.txt",net0.n_2_3_1.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_2_LOCAL.txt",net0.n_2_3_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_2_LOCAL.txt",net0.n_2_3_2.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_2_XPOS.txt",net0.n_2_3_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_2_XNEG.txt",net0.n_2_3_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_2_YPOS.txt",net0.n_2_3_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_2_YNEG.txt",net0.n_2_3_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_2_ZPOS.txt",net0.n_2_3_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_2_ZNEG.txt",net0.n_2_3_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_2_LOCAL.txt",net0.n_2_3_2.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_2_XPOS.txt",net0.n_2_3_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_2_XNEG.txt",net0.n_2_3_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_2_YPOS.txt",net0.n_2_3_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_2_YNEG.txt",net0.n_2_3_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_2_ZPOS.txt",net0.n_2_3_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_2_ZNEG.txt",net0.n_2_3_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_2_LOCAL.txt",net0.n_2_3_2.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_2_XPOS.txt",net0.n_2_3_2.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_2_XNEG.txt",net0.n_2_3_2.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_2_YPOS.txt",net0.n_2_3_2.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_2_YNEG.txt",net0.n_2_3_2.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_2_ZPOS.txt",net0.n_2_3_2.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_2_ZNEG.txt",net0.n_2_3_2.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_2_3_2.txt",net0.n_2_3_2.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_3_LOCAL.txt",net0.n_2_3_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_3_LOCAL.txt",net0.n_2_3_3.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_3_XPOS.txt",net0.n_2_3_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_3_XNEG.txt",net0.n_2_3_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_3_YPOS.txt",net0.n_2_3_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_3_YNEG.txt",net0.n_2_3_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_3_ZPOS.txt",net0.n_2_3_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_2_3_3_ZNEG.txt",net0.n_2_3_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_3_LOCAL.txt",net0.n_2_3_3.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_3_XPOS.txt",net0.n_2_3_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_3_XNEG.txt",net0.n_2_3_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_3_YPOS.txt",net0.n_2_3_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_3_YNEG.txt",net0.n_2_3_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_3_ZPOS.txt",net0.n_2_3_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_2_3_3_ZNEG.txt",net0.n_2_3_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_3_LOCAL.txt",net0.n_2_3_3.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_3_XPOS.txt",net0.n_2_3_3.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_3_XNEG.txt",net0.n_2_3_3.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_3_YPOS.txt",net0.n_2_3_3.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_3_YNEG.txt",net0.n_2_3_3.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_3_ZPOS.txt",net0.n_2_3_3.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_2_3_3_ZNEG.txt",net0.n_2_3_3.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_2_3_3.txt",net0.n_2_3_3.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_0_LOCAL.txt",net0.n_3_0_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_0_LOCAL.txt",net0.n_3_0_0.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_0_XPOS.txt",net0.n_3_0_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_0_XNEG.txt",net0.n_3_0_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_0_YPOS.txt",net0.n_3_0_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_0_YNEG.txt",net0.n_3_0_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_0_ZPOS.txt",net0.n_3_0_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_0_ZNEG.txt",net0.n_3_0_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_0_LOCAL.txt",net0.n_3_0_0.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_0_XPOS.txt",net0.n_3_0_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_0_XNEG.txt",net0.n_3_0_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_0_YPOS.txt",net0.n_3_0_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_0_YNEG.txt",net0.n_3_0_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_0_ZPOS.txt",net0.n_3_0_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_0_ZNEG.txt",net0.n_3_0_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_0_LOCAL.txt",net0.n_3_0_0.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_0_XPOS.txt",net0.n_3_0_0.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_0_XNEG.txt",net0.n_3_0_0.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_0_YPOS.txt",net0.n_3_0_0.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_0_YNEG.txt",net0.n_3_0_0.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_0_ZPOS.txt",net0.n_3_0_0.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_0_ZNEG.txt",net0.n_3_0_0.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_3_0_0.txt",net0.n_3_0_0.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_1_LOCAL.txt",net0.n_3_0_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_1_LOCAL.txt",net0.n_3_0_1.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_1_XPOS.txt",net0.n_3_0_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_1_XNEG.txt",net0.n_3_0_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_1_YPOS.txt",net0.n_3_0_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_1_YNEG.txt",net0.n_3_0_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_1_ZPOS.txt",net0.n_3_0_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_1_ZNEG.txt",net0.n_3_0_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_1_LOCAL.txt",net0.n_3_0_1.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_1_XPOS.txt",net0.n_3_0_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_1_XNEG.txt",net0.n_3_0_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_1_YPOS.txt",net0.n_3_0_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_1_YNEG.txt",net0.n_3_0_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_1_ZPOS.txt",net0.n_3_0_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_1_ZNEG.txt",net0.n_3_0_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_1_LOCAL.txt",net0.n_3_0_1.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_1_XPOS.txt",net0.n_3_0_1.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_1_XNEG.txt",net0.n_3_0_1.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_1_YPOS.txt",net0.n_3_0_1.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_1_YNEG.txt",net0.n_3_0_1.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_1_ZPOS.txt",net0.n_3_0_1.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_1_ZNEG.txt",net0.n_3_0_1.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_3_0_1.txt",net0.n_3_0_1.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_2_LOCAL.txt",net0.n_3_0_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_2_LOCAL.txt",net0.n_3_0_2.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_2_XPOS.txt",net0.n_3_0_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_2_XNEG.txt",net0.n_3_0_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_2_YPOS.txt",net0.n_3_0_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_2_YNEG.txt",net0.n_3_0_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_2_ZPOS.txt",net0.n_3_0_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_2_ZNEG.txt",net0.n_3_0_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_2_LOCAL.txt",net0.n_3_0_2.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_2_XPOS.txt",net0.n_3_0_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_2_XNEG.txt",net0.n_3_0_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_2_YPOS.txt",net0.n_3_0_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_2_YNEG.txt",net0.n_3_0_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_2_ZPOS.txt",net0.n_3_0_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_2_ZNEG.txt",net0.n_3_0_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_2_LOCAL.txt",net0.n_3_0_2.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_2_XPOS.txt",net0.n_3_0_2.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_2_XNEG.txt",net0.n_3_0_2.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_2_YPOS.txt",net0.n_3_0_2.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_2_YNEG.txt",net0.n_3_0_2.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_2_ZPOS.txt",net0.n_3_0_2.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_2_ZNEG.txt",net0.n_3_0_2.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_3_0_2.txt",net0.n_3_0_2.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_3_LOCAL.txt",net0.n_3_0_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_3_LOCAL.txt",net0.n_3_0_3.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_3_XPOS.txt",net0.n_3_0_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_3_XNEG.txt",net0.n_3_0_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_3_YPOS.txt",net0.n_3_0_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_3_YNEG.txt",net0.n_3_0_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_3_ZPOS.txt",net0.n_3_0_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_0_3_ZNEG.txt",net0.n_3_0_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_3_LOCAL.txt",net0.n_3_0_3.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_3_XPOS.txt",net0.n_3_0_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_3_XNEG.txt",net0.n_3_0_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_3_YPOS.txt",net0.n_3_0_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_3_YNEG.txt",net0.n_3_0_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_3_ZPOS.txt",net0.n_3_0_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_0_3_ZNEG.txt",net0.n_3_0_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_3_LOCAL.txt",net0.n_3_0_3.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_3_XPOS.txt",net0.n_3_0_3.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_3_XNEG.txt",net0.n_3_0_3.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_3_YPOS.txt",net0.n_3_0_3.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_3_YNEG.txt",net0.n_3_0_3.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_3_ZPOS.txt",net0.n_3_0_3.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_0_3_ZNEG.txt",net0.n_3_0_3.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_3_0_3.txt",net0.n_3_0_3.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_0_LOCAL.txt",net0.n_3_1_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_0_LOCAL.txt",net0.n_3_1_0.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_0_XPOS.txt",net0.n_3_1_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_0_XNEG.txt",net0.n_3_1_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_0_YPOS.txt",net0.n_3_1_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_0_YNEG.txt",net0.n_3_1_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_0_ZPOS.txt",net0.n_3_1_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_0_ZNEG.txt",net0.n_3_1_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_0_LOCAL.txt",net0.n_3_1_0.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_0_XPOS.txt",net0.n_3_1_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_0_XNEG.txt",net0.n_3_1_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_0_YPOS.txt",net0.n_3_1_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_0_YNEG.txt",net0.n_3_1_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_0_ZPOS.txt",net0.n_3_1_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_0_ZNEG.txt",net0.n_3_1_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_0_LOCAL.txt",net0.n_3_1_0.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_0_XPOS.txt",net0.n_3_1_0.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_0_XNEG.txt",net0.n_3_1_0.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_0_YPOS.txt",net0.n_3_1_0.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_0_YNEG.txt",net0.n_3_1_0.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_0_ZPOS.txt",net0.n_3_1_0.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_0_ZNEG.txt",net0.n_3_1_0.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_3_1_0.txt",net0.n_3_1_0.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_1_LOCAL.txt",net0.n_3_1_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_1_LOCAL.txt",net0.n_3_1_1.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_1_XPOS.txt",net0.n_3_1_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_1_XNEG.txt",net0.n_3_1_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_1_YPOS.txt",net0.n_3_1_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_1_YNEG.txt",net0.n_3_1_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_1_ZPOS.txt",net0.n_3_1_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_1_ZNEG.txt",net0.n_3_1_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_1_LOCAL.txt",net0.n_3_1_1.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_1_XPOS.txt",net0.n_3_1_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_1_XNEG.txt",net0.n_3_1_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_1_YPOS.txt",net0.n_3_1_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_1_YNEG.txt",net0.n_3_1_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_1_ZPOS.txt",net0.n_3_1_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_1_ZNEG.txt",net0.n_3_1_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_1_LOCAL.txt",net0.n_3_1_1.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_1_XPOS.txt",net0.n_3_1_1.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_1_XNEG.txt",net0.n_3_1_1.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_1_YPOS.txt",net0.n_3_1_1.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_1_YNEG.txt",net0.n_3_1_1.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_1_ZPOS.txt",net0.n_3_1_1.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_1_ZNEG.txt",net0.n_3_1_1.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_3_1_1.txt",net0.n_3_1_1.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_2_LOCAL.txt",net0.n_3_1_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_2_LOCAL.txt",net0.n_3_1_2.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_2_XPOS.txt",net0.n_3_1_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_2_XNEG.txt",net0.n_3_1_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_2_YPOS.txt",net0.n_3_1_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_2_YNEG.txt",net0.n_3_1_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_2_ZPOS.txt",net0.n_3_1_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_2_ZNEG.txt",net0.n_3_1_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_2_LOCAL.txt",net0.n_3_1_2.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_2_XPOS.txt",net0.n_3_1_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_2_XNEG.txt",net0.n_3_1_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_2_YPOS.txt",net0.n_3_1_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_2_YNEG.txt",net0.n_3_1_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_2_ZPOS.txt",net0.n_3_1_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_2_ZNEG.txt",net0.n_3_1_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_2_LOCAL.txt",net0.n_3_1_2.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_2_XPOS.txt",net0.n_3_1_2.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_2_XNEG.txt",net0.n_3_1_2.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_2_YPOS.txt",net0.n_3_1_2.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_2_YNEG.txt",net0.n_3_1_2.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_2_ZPOS.txt",net0.n_3_1_2.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_2_ZNEG.txt",net0.n_3_1_2.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_3_1_2.txt",net0.n_3_1_2.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_3_LOCAL.txt",net0.n_3_1_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_3_LOCAL.txt",net0.n_3_1_3.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_3_XPOS.txt",net0.n_3_1_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_3_XNEG.txt",net0.n_3_1_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_3_YPOS.txt",net0.n_3_1_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_3_YNEG.txt",net0.n_3_1_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_3_ZPOS.txt",net0.n_3_1_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_1_3_ZNEG.txt",net0.n_3_1_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_3_LOCAL.txt",net0.n_3_1_3.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_3_XPOS.txt",net0.n_3_1_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_3_XNEG.txt",net0.n_3_1_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_3_YPOS.txt",net0.n_3_1_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_3_YNEG.txt",net0.n_3_1_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_3_ZPOS.txt",net0.n_3_1_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_1_3_ZNEG.txt",net0.n_3_1_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_3_LOCAL.txt",net0.n_3_1_3.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_3_XPOS.txt",net0.n_3_1_3.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_3_XNEG.txt",net0.n_3_1_3.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_3_YPOS.txt",net0.n_3_1_3.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_3_YNEG.txt",net0.n_3_1_3.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_3_ZPOS.txt",net0.n_3_1_3.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_1_3_ZNEG.txt",net0.n_3_1_3.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_3_1_3.txt",net0.n_3_1_3.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_0_LOCAL.txt",net0.n_3_2_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_0_LOCAL.txt",net0.n_3_2_0.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_0_XPOS.txt",net0.n_3_2_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_0_XNEG.txt",net0.n_3_2_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_0_YPOS.txt",net0.n_3_2_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_0_YNEG.txt",net0.n_3_2_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_0_ZPOS.txt",net0.n_3_2_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_0_ZNEG.txt",net0.n_3_2_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_0_LOCAL.txt",net0.n_3_2_0.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_0_XPOS.txt",net0.n_3_2_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_0_XNEG.txt",net0.n_3_2_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_0_YPOS.txt",net0.n_3_2_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_0_YNEG.txt",net0.n_3_2_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_0_ZPOS.txt",net0.n_3_2_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_0_ZNEG.txt",net0.n_3_2_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_0_LOCAL.txt",net0.n_3_2_0.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_0_XPOS.txt",net0.n_3_2_0.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_0_XNEG.txt",net0.n_3_2_0.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_0_YPOS.txt",net0.n_3_2_0.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_0_YNEG.txt",net0.n_3_2_0.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_0_ZPOS.txt",net0.n_3_2_0.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_0_ZNEG.txt",net0.n_3_2_0.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_3_2_0.txt",net0.n_3_2_0.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_1_LOCAL.txt",net0.n_3_2_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_1_LOCAL.txt",net0.n_3_2_1.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_1_XPOS.txt",net0.n_3_2_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_1_XNEG.txt",net0.n_3_2_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_1_YPOS.txt",net0.n_3_2_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_1_YNEG.txt",net0.n_3_2_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_1_ZPOS.txt",net0.n_3_2_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_1_ZNEG.txt",net0.n_3_2_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_1_LOCAL.txt",net0.n_3_2_1.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_1_XPOS.txt",net0.n_3_2_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_1_XNEG.txt",net0.n_3_2_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_1_YPOS.txt",net0.n_3_2_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_1_YNEG.txt",net0.n_3_2_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_1_ZPOS.txt",net0.n_3_2_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_1_ZNEG.txt",net0.n_3_2_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_1_LOCAL.txt",net0.n_3_2_1.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_1_XPOS.txt",net0.n_3_2_1.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_1_XNEG.txt",net0.n_3_2_1.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_1_YPOS.txt",net0.n_3_2_1.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_1_YNEG.txt",net0.n_3_2_1.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_1_ZPOS.txt",net0.n_3_2_1.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_1_ZNEG.txt",net0.n_3_2_1.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_3_2_1.txt",net0.n_3_2_1.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_2_LOCAL.txt",net0.n_3_2_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_2_LOCAL.txt",net0.n_3_2_2.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_2_XPOS.txt",net0.n_3_2_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_2_XNEG.txt",net0.n_3_2_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_2_YPOS.txt",net0.n_3_2_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_2_YNEG.txt",net0.n_3_2_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_2_ZPOS.txt",net0.n_3_2_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_2_ZNEG.txt",net0.n_3_2_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_2_LOCAL.txt",net0.n_3_2_2.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_2_XPOS.txt",net0.n_3_2_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_2_XNEG.txt",net0.n_3_2_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_2_YPOS.txt",net0.n_3_2_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_2_YNEG.txt",net0.n_3_2_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_2_ZPOS.txt",net0.n_3_2_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_2_ZNEG.txt",net0.n_3_2_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_2_LOCAL.txt",net0.n_3_2_2.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_2_XPOS.txt",net0.n_3_2_2.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_2_XNEG.txt",net0.n_3_2_2.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_2_YPOS.txt",net0.n_3_2_2.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_2_YNEG.txt",net0.n_3_2_2.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_2_ZPOS.txt",net0.n_3_2_2.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_2_ZNEG.txt",net0.n_3_2_2.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_3_2_2.txt",net0.n_3_2_2.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_3_LOCAL.txt",net0.n_3_2_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_3_LOCAL.txt",net0.n_3_2_3.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_3_XPOS.txt",net0.n_3_2_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_3_XNEG.txt",net0.n_3_2_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_3_YPOS.txt",net0.n_3_2_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_3_YNEG.txt",net0.n_3_2_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_3_ZPOS.txt",net0.n_3_2_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_2_3_ZNEG.txt",net0.n_3_2_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_3_LOCAL.txt",net0.n_3_2_3.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_3_XPOS.txt",net0.n_3_2_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_3_XNEG.txt",net0.n_3_2_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_3_YPOS.txt",net0.n_3_2_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_3_YNEG.txt",net0.n_3_2_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_3_ZPOS.txt",net0.n_3_2_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_2_3_ZNEG.txt",net0.n_3_2_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_3_LOCAL.txt",net0.n_3_2_3.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_3_XPOS.txt",net0.n_3_2_3.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_3_XNEG.txt",net0.n_3_2_3.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_3_YPOS.txt",net0.n_3_2_3.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_3_YNEG.txt",net0.n_3_2_3.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_3_ZPOS.txt",net0.n_3_2_3.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_2_3_ZNEG.txt",net0.n_3_2_3.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_3_2_3.txt",net0.n_3_2_3.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_0_LOCAL.txt",net0.n_3_3_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_0_LOCAL.txt",net0.n_3_3_0.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_0_XPOS.txt",net0.n_3_3_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_0_XNEG.txt",net0.n_3_3_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_0_YPOS.txt",net0.n_3_3_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_0_YNEG.txt",net0.n_3_3_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_0_ZPOS.txt",net0.n_3_3_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_0_ZNEG.txt",net0.n_3_3_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_0_LOCAL.txt",net0.n_3_3_0.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_0_XPOS.txt",net0.n_3_3_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_0_XNEG.txt",net0.n_3_3_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_0_YPOS.txt",net0.n_3_3_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_0_YNEG.txt",net0.n_3_3_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_0_ZPOS.txt",net0.n_3_3_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_0_ZNEG.txt",net0.n_3_3_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_0_LOCAL.txt",net0.n_3_3_0.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_0_XPOS.txt",net0.n_3_3_0.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_0_XNEG.txt",net0.n_3_3_0.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_0_YPOS.txt",net0.n_3_3_0.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_0_YNEG.txt",net0.n_3_3_0.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_0_ZPOS.txt",net0.n_3_3_0.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_0_ZNEG.txt",net0.n_3_3_0.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_3_3_0.txt",net0.n_3_3_0.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_1_LOCAL.txt",net0.n_3_3_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_1_LOCAL.txt",net0.n_3_3_1.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_1_XPOS.txt",net0.n_3_3_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_1_XNEG.txt",net0.n_3_3_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_1_YPOS.txt",net0.n_3_3_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_1_YNEG.txt",net0.n_3_3_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_1_ZPOS.txt",net0.n_3_3_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_1_ZNEG.txt",net0.n_3_3_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_1_LOCAL.txt",net0.n_3_3_1.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_1_XPOS.txt",net0.n_3_3_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_1_XNEG.txt",net0.n_3_3_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_1_YPOS.txt",net0.n_3_3_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_1_YNEG.txt",net0.n_3_3_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_1_ZPOS.txt",net0.n_3_3_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_1_ZNEG.txt",net0.n_3_3_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_1_LOCAL.txt",net0.n_3_3_1.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_1_XPOS.txt",net0.n_3_3_1.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_1_XNEG.txt",net0.n_3_3_1.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_1_YPOS.txt",net0.n_3_3_1.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_1_YNEG.txt",net0.n_3_3_1.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_1_ZPOS.txt",net0.n_3_3_1.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_1_ZNEG.txt",net0.n_3_3_1.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_3_3_1.txt",net0.n_3_3_1.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_2_LOCAL.txt",net0.n_3_3_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_2_LOCAL.txt",net0.n_3_3_2.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_2_XPOS.txt",net0.n_3_3_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_2_XNEG.txt",net0.n_3_3_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_2_YPOS.txt",net0.n_3_3_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_2_YNEG.txt",net0.n_3_3_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_2_ZPOS.txt",net0.n_3_3_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_2_ZNEG.txt",net0.n_3_3_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_2_LOCAL.txt",net0.n_3_3_2.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_2_XPOS.txt",net0.n_3_3_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_2_XNEG.txt",net0.n_3_3_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_2_YPOS.txt",net0.n_3_3_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_2_YNEG.txt",net0.n_3_3_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_2_ZPOS.txt",net0.n_3_3_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_2_ZNEG.txt",net0.n_3_3_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_2_LOCAL.txt",net0.n_3_3_2.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_2_XPOS.txt",net0.n_3_3_2.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_2_XNEG.txt",net0.n_3_3_2.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_2_YPOS.txt",net0.n_3_3_2.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_2_YNEG.txt",net0.n_3_3_2.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_2_ZPOS.txt",net0.n_3_3_2.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_2_ZNEG.txt",net0.n_3_3_2.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_3_3_2.txt",net0.n_3_3_2.local_unit_inst.data);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_3_LOCAL.txt",net0.n_3_3_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_3_LOCAL.txt",net0.n_3_3_3.switch_inst.LOCAL.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_3_XPOS.txt",net0.n_3_3_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_3_XNEG.txt",net0.n_3_3_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_3_YPOS.txt",net0.n_3_3_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_3_YNEG.txt",net0.n_3_3_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_3_ZPOS.txt",net0.n_3_3_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/routing_table_3_3_3_ZNEG.txt",net0.n_3_3_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_3_LOCAL.txt",net0.n_3_3_3.switch_inst.LOCAL.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_3_XPOS.txt",net0.n_3_3_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_3_XNEG.txt",net0.n_3_3_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_3_YPOS.txt",net0.n_3_3_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_3_YNEG.txt",net0.n_3_3_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_3_ZPOS.txt",net0.n_3_3_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/multicast_table_3_3_3_ZNEG.txt",net0.n_3_3_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_3_LOCAL.txt",net0.n_3_3_3.switch_inst.mux_local.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_3_XPOS.txt",net0.n_3_3_3.switch_inst.mux_xpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_3_XNEG.txt",net0.n_3_3_3.switch_inst.mux_xneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_3_YPOS.txt",net0.n_3_3_3.switch_inst.mux_ypos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_3_YNEG.txt",net0.n_3_3_3.switch_inst.mux_yneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_3_ZPOS.txt",net0.n_3_3_3.switch_inst.mux_zpos.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/tables/reduction_table_3_3_3_ZNEG.txt",net0.n_3_3_3.switch_inst.mux_zneg.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction_data/input_data/data_to_send_3_3_3.txt",net0.n_3_3_3.local_unit_inst.data);
	initial begin
		clk=0;
		rst=1;

		#100 rst=0;
	end
endmodule
