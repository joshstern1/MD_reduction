module network_tb;
	parameter PayloadLen=128;
    parameter DataWidth=256;
    parameter WeightPos=144;
    parameter WeightWidth=8;
    parameter IndexPos=128;
    parameter IndexWidth=16;
    parameter PriorityPos=152;
    parameter PriorityWidth=8;
    parameter ExitPos=160;
    parameter ExitWidth=4;
    parameter InterNodeFIFODepth=128;
    parameter IntraNodeFIFODepth=1;
    parameter RoutingTableWidth=32;
    parameter RoutingTablesize=256;
    parameter MulticastTableWidth=103;
    parameter MulticastTablesize=256;
    parameter ReductionTableWidth=162;
    parameter ReductionTablesize=256;
    parameter PcktTypeLen=4;
    parameter profiling_freq=10;


 	reg clk,rst;

	always #5 clk=~clk;

	network net0(clk,rst);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_0_local.txt",net0.n_0_0_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_0_xpos.txt",net0.n_0_0_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_0_xneg.txt",net0.n_0_0_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_0_ypos.txt",net0.n_0_0_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_0_yneg.txt",net0.n_0_0_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_0_zpos.txt",net0.n_0_0_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_0_zneg.txt",net0.n_0_0_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_0_xpos.txt",net0.n_0_0_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_0_xneg.txt",net0.n_0_0_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_0_ypos.txt",net0.n_0_0_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_0_yneg.txt",net0.n_0_0_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_0_zpos.txt",net0.n_0_0_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_0_zneg.txt",net0.n_0_0_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_0_xpos.txt",net0.n_0_0_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_0_xneg.txt",net0.n_0_0_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_0_ypos.txt",net0.n_0_0_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_0_yneg.txt",net0.n_0_0_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_0_zpos.txt",net0.n_0_0_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_0_zneg.txt",net0.n_0_0_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_1_local.txt",net0.n_0_0_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_1_xpos.txt",net0.n_0_0_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_1_xneg.txt",net0.n_0_0_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_1_ypos.txt",net0.n_0_0_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_1_yneg.txt",net0.n_0_0_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_1_zpos.txt",net0.n_0_0_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_1_zneg.txt",net0.n_0_0_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_1_xpos.txt",net0.n_0_0_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_1_xneg.txt",net0.n_0_0_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_1_ypos.txt",net0.n_0_0_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_1_yneg.txt",net0.n_0_0_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_1_zpos.txt",net0.n_0_0_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_1_zneg.txt",net0.n_0_0_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_1_xpos.txt",net0.n_0_0_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_1_xneg.txt",net0.n_0_0_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_1_ypos.txt",net0.n_0_0_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_1_yneg.txt",net0.n_0_0_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_1_zpos.txt",net0.n_0_0_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_1_zneg.txt",net0.n_0_0_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_2_local.txt",net0.n_0_0_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_2_xpos.txt",net0.n_0_0_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_2_xneg.txt",net0.n_0_0_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_2_ypos.txt",net0.n_0_0_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_2_yneg.txt",net0.n_0_0_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_2_zpos.txt",net0.n_0_0_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_2_zneg.txt",net0.n_0_0_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_2_xpos.txt",net0.n_0_0_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_2_xneg.txt",net0.n_0_0_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_2_ypos.txt",net0.n_0_0_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_2_yneg.txt",net0.n_0_0_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_2_zpos.txt",net0.n_0_0_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_2_zneg.txt",net0.n_0_0_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_2_xpos.txt",net0.n_0_0_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_2_xneg.txt",net0.n_0_0_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_2_ypos.txt",net0.n_0_0_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_2_yneg.txt",net0.n_0_0_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_2_zpos.txt",net0.n_0_0_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_2_zneg.txt",net0.n_0_0_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_3_local.txt",net0.n_0_0_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_3_xpos.txt",net0.n_0_0_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_3_xneg.txt",net0.n_0_0_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_3_ypos.txt",net0.n_0_0_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_3_yneg.txt",net0.n_0_0_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_3_zpos.txt",net0.n_0_0_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_3_zneg.txt",net0.n_0_0_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_3_xpos.txt",net0.n_0_0_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_3_xneg.txt",net0.n_0_0_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_3_ypos.txt",net0.n_0_0_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_3_yneg.txt",net0.n_0_0_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_3_zpos.txt",net0.n_0_0_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_3_zneg.txt",net0.n_0_0_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_3_xpos.txt",net0.n_0_0_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_3_xneg.txt",net0.n_0_0_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_3_ypos.txt",net0.n_0_0_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_3_yneg.txt",net0.n_0_0_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_3_zpos.txt",net0.n_0_0_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_3_zneg.txt",net0.n_0_0_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_4_local.txt",net0.n_0_0_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_4_xpos.txt",net0.n_0_0_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_4_xneg.txt",net0.n_0_0_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_4_ypos.txt",net0.n_0_0_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_4_yneg.txt",net0.n_0_0_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_4_zpos.txt",net0.n_0_0_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_4_zneg.txt",net0.n_0_0_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_4_xpos.txt",net0.n_0_0_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_4_xneg.txt",net0.n_0_0_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_4_ypos.txt",net0.n_0_0_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_4_yneg.txt",net0.n_0_0_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_4_zpos.txt",net0.n_0_0_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_4_zneg.txt",net0.n_0_0_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_4_xpos.txt",net0.n_0_0_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_4_xneg.txt",net0.n_0_0_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_4_ypos.txt",net0.n_0_0_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_4_yneg.txt",net0.n_0_0_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_4_zpos.txt",net0.n_0_0_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_4_zneg.txt",net0.n_0_0_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_5_local.txt",net0.n_0_0_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_5_xpos.txt",net0.n_0_0_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_5_xneg.txt",net0.n_0_0_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_5_ypos.txt",net0.n_0_0_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_5_yneg.txt",net0.n_0_0_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_5_zpos.txt",net0.n_0_0_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_5_zneg.txt",net0.n_0_0_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_5_xpos.txt",net0.n_0_0_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_5_xneg.txt",net0.n_0_0_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_5_ypos.txt",net0.n_0_0_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_5_yneg.txt",net0.n_0_0_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_5_zpos.txt",net0.n_0_0_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_5_zneg.txt",net0.n_0_0_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_5_xpos.txt",net0.n_0_0_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_5_xneg.txt",net0.n_0_0_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_5_ypos.txt",net0.n_0_0_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_5_yneg.txt",net0.n_0_0_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_5_zpos.txt",net0.n_0_0_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_5_zneg.txt",net0.n_0_0_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_6_local.txt",net0.n_0_0_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_6_xpos.txt",net0.n_0_0_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_6_xneg.txt",net0.n_0_0_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_6_ypos.txt",net0.n_0_0_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_6_yneg.txt",net0.n_0_0_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_6_zpos.txt",net0.n_0_0_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_6_zneg.txt",net0.n_0_0_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_6_xpos.txt",net0.n_0_0_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_6_xneg.txt",net0.n_0_0_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_6_ypos.txt",net0.n_0_0_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_6_yneg.txt",net0.n_0_0_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_6_zpos.txt",net0.n_0_0_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_6_zneg.txt",net0.n_0_0_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_6_xpos.txt",net0.n_0_0_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_6_xneg.txt",net0.n_0_0_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_6_ypos.txt",net0.n_0_0_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_6_yneg.txt",net0.n_0_0_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_6_zpos.txt",net0.n_0_0_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_6_zneg.txt",net0.n_0_0_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_7_local.txt",net0.n_0_0_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_7_xpos.txt",net0.n_0_0_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_7_xneg.txt",net0.n_0_0_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_7_ypos.txt",net0.n_0_0_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_7_yneg.txt",net0.n_0_0_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_7_zpos.txt",net0.n_0_0_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_0_7_zneg.txt",net0.n_0_0_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_7_xpos.txt",net0.n_0_0_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_7_xneg.txt",net0.n_0_0_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_7_ypos.txt",net0.n_0_0_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_7_yneg.txt",net0.n_0_0_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_7_zpos.txt",net0.n_0_0_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_0_7_zneg.txt",net0.n_0_0_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_7_xpos.txt",net0.n_0_0_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_7_xneg.txt",net0.n_0_0_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_7_ypos.txt",net0.n_0_0_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_7_yneg.txt",net0.n_0_0_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_7_zpos.txt",net0.n_0_0_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_0_7_zneg.txt",net0.n_0_0_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_0_local.txt",net0.n_0_1_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_0_xpos.txt",net0.n_0_1_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_0_xneg.txt",net0.n_0_1_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_0_ypos.txt",net0.n_0_1_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_0_yneg.txt",net0.n_0_1_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_0_zpos.txt",net0.n_0_1_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_0_zneg.txt",net0.n_0_1_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_0_xpos.txt",net0.n_0_1_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_0_xneg.txt",net0.n_0_1_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_0_ypos.txt",net0.n_0_1_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_0_yneg.txt",net0.n_0_1_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_0_zpos.txt",net0.n_0_1_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_0_zneg.txt",net0.n_0_1_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_0_xpos.txt",net0.n_0_1_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_0_xneg.txt",net0.n_0_1_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_0_ypos.txt",net0.n_0_1_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_0_yneg.txt",net0.n_0_1_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_0_zpos.txt",net0.n_0_1_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_0_zneg.txt",net0.n_0_1_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_1_local.txt",net0.n_0_1_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_1_xpos.txt",net0.n_0_1_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_1_xneg.txt",net0.n_0_1_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_1_ypos.txt",net0.n_0_1_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_1_yneg.txt",net0.n_0_1_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_1_zpos.txt",net0.n_0_1_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_1_zneg.txt",net0.n_0_1_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_1_xpos.txt",net0.n_0_1_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_1_xneg.txt",net0.n_0_1_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_1_ypos.txt",net0.n_0_1_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_1_yneg.txt",net0.n_0_1_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_1_zpos.txt",net0.n_0_1_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_1_zneg.txt",net0.n_0_1_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_1_xpos.txt",net0.n_0_1_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_1_xneg.txt",net0.n_0_1_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_1_ypos.txt",net0.n_0_1_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_1_yneg.txt",net0.n_0_1_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_1_zpos.txt",net0.n_0_1_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_1_zneg.txt",net0.n_0_1_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_2_local.txt",net0.n_0_1_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_2_xpos.txt",net0.n_0_1_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_2_xneg.txt",net0.n_0_1_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_2_ypos.txt",net0.n_0_1_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_2_yneg.txt",net0.n_0_1_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_2_zpos.txt",net0.n_0_1_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_2_zneg.txt",net0.n_0_1_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_2_xpos.txt",net0.n_0_1_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_2_xneg.txt",net0.n_0_1_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_2_ypos.txt",net0.n_0_1_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_2_yneg.txt",net0.n_0_1_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_2_zpos.txt",net0.n_0_1_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_2_zneg.txt",net0.n_0_1_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_2_xpos.txt",net0.n_0_1_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_2_xneg.txt",net0.n_0_1_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_2_ypos.txt",net0.n_0_1_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_2_yneg.txt",net0.n_0_1_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_2_zpos.txt",net0.n_0_1_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_2_zneg.txt",net0.n_0_1_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_3_local.txt",net0.n_0_1_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_3_xpos.txt",net0.n_0_1_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_3_xneg.txt",net0.n_0_1_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_3_ypos.txt",net0.n_0_1_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_3_yneg.txt",net0.n_0_1_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_3_zpos.txt",net0.n_0_1_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_3_zneg.txt",net0.n_0_1_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_3_xpos.txt",net0.n_0_1_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_3_xneg.txt",net0.n_0_1_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_3_ypos.txt",net0.n_0_1_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_3_yneg.txt",net0.n_0_1_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_3_zpos.txt",net0.n_0_1_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_3_zneg.txt",net0.n_0_1_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_3_xpos.txt",net0.n_0_1_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_3_xneg.txt",net0.n_0_1_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_3_ypos.txt",net0.n_0_1_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_3_yneg.txt",net0.n_0_1_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_3_zpos.txt",net0.n_0_1_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_3_zneg.txt",net0.n_0_1_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_4_local.txt",net0.n_0_1_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_4_xpos.txt",net0.n_0_1_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_4_xneg.txt",net0.n_0_1_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_4_ypos.txt",net0.n_0_1_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_4_yneg.txt",net0.n_0_1_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_4_zpos.txt",net0.n_0_1_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_4_zneg.txt",net0.n_0_1_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_4_xpos.txt",net0.n_0_1_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_4_xneg.txt",net0.n_0_1_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_4_ypos.txt",net0.n_0_1_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_4_yneg.txt",net0.n_0_1_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_4_zpos.txt",net0.n_0_1_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_4_zneg.txt",net0.n_0_1_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_4_xpos.txt",net0.n_0_1_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_4_xneg.txt",net0.n_0_1_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_4_ypos.txt",net0.n_0_1_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_4_yneg.txt",net0.n_0_1_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_4_zpos.txt",net0.n_0_1_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_4_zneg.txt",net0.n_0_1_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_5_local.txt",net0.n_0_1_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_5_xpos.txt",net0.n_0_1_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_5_xneg.txt",net0.n_0_1_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_5_ypos.txt",net0.n_0_1_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_5_yneg.txt",net0.n_0_1_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_5_zpos.txt",net0.n_0_1_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_5_zneg.txt",net0.n_0_1_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_5_xpos.txt",net0.n_0_1_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_5_xneg.txt",net0.n_0_1_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_5_ypos.txt",net0.n_0_1_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_5_yneg.txt",net0.n_0_1_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_5_zpos.txt",net0.n_0_1_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_5_zneg.txt",net0.n_0_1_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_5_xpos.txt",net0.n_0_1_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_5_xneg.txt",net0.n_0_1_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_5_ypos.txt",net0.n_0_1_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_5_yneg.txt",net0.n_0_1_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_5_zpos.txt",net0.n_0_1_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_5_zneg.txt",net0.n_0_1_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_6_local.txt",net0.n_0_1_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_6_xpos.txt",net0.n_0_1_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_6_xneg.txt",net0.n_0_1_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_6_ypos.txt",net0.n_0_1_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_6_yneg.txt",net0.n_0_1_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_6_zpos.txt",net0.n_0_1_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_6_zneg.txt",net0.n_0_1_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_6_xpos.txt",net0.n_0_1_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_6_xneg.txt",net0.n_0_1_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_6_ypos.txt",net0.n_0_1_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_6_yneg.txt",net0.n_0_1_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_6_zpos.txt",net0.n_0_1_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_6_zneg.txt",net0.n_0_1_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_6_xpos.txt",net0.n_0_1_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_6_xneg.txt",net0.n_0_1_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_6_ypos.txt",net0.n_0_1_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_6_yneg.txt",net0.n_0_1_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_6_zpos.txt",net0.n_0_1_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_6_zneg.txt",net0.n_0_1_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_7_local.txt",net0.n_0_1_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_7_xpos.txt",net0.n_0_1_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_7_xneg.txt",net0.n_0_1_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_7_ypos.txt",net0.n_0_1_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_7_yneg.txt",net0.n_0_1_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_7_zpos.txt",net0.n_0_1_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_1_7_zneg.txt",net0.n_0_1_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_7_xpos.txt",net0.n_0_1_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_7_xneg.txt",net0.n_0_1_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_7_ypos.txt",net0.n_0_1_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_7_yneg.txt",net0.n_0_1_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_7_zpos.txt",net0.n_0_1_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_1_7_zneg.txt",net0.n_0_1_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_7_xpos.txt",net0.n_0_1_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_7_xneg.txt",net0.n_0_1_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_7_ypos.txt",net0.n_0_1_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_7_yneg.txt",net0.n_0_1_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_7_zpos.txt",net0.n_0_1_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_1_7_zneg.txt",net0.n_0_1_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_0_local.txt",net0.n_0_2_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_0_xpos.txt",net0.n_0_2_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_0_xneg.txt",net0.n_0_2_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_0_ypos.txt",net0.n_0_2_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_0_yneg.txt",net0.n_0_2_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_0_zpos.txt",net0.n_0_2_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_0_zneg.txt",net0.n_0_2_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_0_xpos.txt",net0.n_0_2_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_0_xneg.txt",net0.n_0_2_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_0_ypos.txt",net0.n_0_2_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_0_yneg.txt",net0.n_0_2_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_0_zpos.txt",net0.n_0_2_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_0_zneg.txt",net0.n_0_2_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_0_xpos.txt",net0.n_0_2_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_0_xneg.txt",net0.n_0_2_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_0_ypos.txt",net0.n_0_2_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_0_yneg.txt",net0.n_0_2_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_0_zpos.txt",net0.n_0_2_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_0_zneg.txt",net0.n_0_2_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_1_local.txt",net0.n_0_2_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_1_xpos.txt",net0.n_0_2_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_1_xneg.txt",net0.n_0_2_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_1_ypos.txt",net0.n_0_2_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_1_yneg.txt",net0.n_0_2_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_1_zpos.txt",net0.n_0_2_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_1_zneg.txt",net0.n_0_2_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_1_xpos.txt",net0.n_0_2_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_1_xneg.txt",net0.n_0_2_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_1_ypos.txt",net0.n_0_2_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_1_yneg.txt",net0.n_0_2_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_1_zpos.txt",net0.n_0_2_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_1_zneg.txt",net0.n_0_2_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_1_xpos.txt",net0.n_0_2_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_1_xneg.txt",net0.n_0_2_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_1_ypos.txt",net0.n_0_2_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_1_yneg.txt",net0.n_0_2_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_1_zpos.txt",net0.n_0_2_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_1_zneg.txt",net0.n_0_2_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_2_local.txt",net0.n_0_2_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_2_xpos.txt",net0.n_0_2_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_2_xneg.txt",net0.n_0_2_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_2_ypos.txt",net0.n_0_2_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_2_yneg.txt",net0.n_0_2_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_2_zpos.txt",net0.n_0_2_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_2_zneg.txt",net0.n_0_2_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_2_xpos.txt",net0.n_0_2_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_2_xneg.txt",net0.n_0_2_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_2_ypos.txt",net0.n_0_2_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_2_yneg.txt",net0.n_0_2_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_2_zpos.txt",net0.n_0_2_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_2_zneg.txt",net0.n_0_2_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_2_xpos.txt",net0.n_0_2_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_2_xneg.txt",net0.n_0_2_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_2_ypos.txt",net0.n_0_2_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_2_yneg.txt",net0.n_0_2_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_2_zpos.txt",net0.n_0_2_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_2_zneg.txt",net0.n_0_2_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_3_local.txt",net0.n_0_2_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_3_xpos.txt",net0.n_0_2_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_3_xneg.txt",net0.n_0_2_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_3_ypos.txt",net0.n_0_2_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_3_yneg.txt",net0.n_0_2_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_3_zpos.txt",net0.n_0_2_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_3_zneg.txt",net0.n_0_2_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_3_xpos.txt",net0.n_0_2_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_3_xneg.txt",net0.n_0_2_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_3_ypos.txt",net0.n_0_2_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_3_yneg.txt",net0.n_0_2_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_3_zpos.txt",net0.n_0_2_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_3_zneg.txt",net0.n_0_2_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_3_xpos.txt",net0.n_0_2_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_3_xneg.txt",net0.n_0_2_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_3_ypos.txt",net0.n_0_2_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_3_yneg.txt",net0.n_0_2_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_3_zpos.txt",net0.n_0_2_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_3_zneg.txt",net0.n_0_2_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_4_local.txt",net0.n_0_2_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_4_xpos.txt",net0.n_0_2_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_4_xneg.txt",net0.n_0_2_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_4_ypos.txt",net0.n_0_2_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_4_yneg.txt",net0.n_0_2_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_4_zpos.txt",net0.n_0_2_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_4_zneg.txt",net0.n_0_2_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_4_xpos.txt",net0.n_0_2_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_4_xneg.txt",net0.n_0_2_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_4_ypos.txt",net0.n_0_2_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_4_yneg.txt",net0.n_0_2_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_4_zpos.txt",net0.n_0_2_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_4_zneg.txt",net0.n_0_2_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_4_xpos.txt",net0.n_0_2_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_4_xneg.txt",net0.n_0_2_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_4_ypos.txt",net0.n_0_2_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_4_yneg.txt",net0.n_0_2_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_4_zpos.txt",net0.n_0_2_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_4_zneg.txt",net0.n_0_2_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_5_local.txt",net0.n_0_2_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_5_xpos.txt",net0.n_0_2_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_5_xneg.txt",net0.n_0_2_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_5_ypos.txt",net0.n_0_2_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_5_yneg.txt",net0.n_0_2_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_5_zpos.txt",net0.n_0_2_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_5_zneg.txt",net0.n_0_2_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_5_xpos.txt",net0.n_0_2_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_5_xneg.txt",net0.n_0_2_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_5_ypos.txt",net0.n_0_2_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_5_yneg.txt",net0.n_0_2_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_5_zpos.txt",net0.n_0_2_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_5_zneg.txt",net0.n_0_2_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_5_xpos.txt",net0.n_0_2_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_5_xneg.txt",net0.n_0_2_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_5_ypos.txt",net0.n_0_2_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_5_yneg.txt",net0.n_0_2_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_5_zpos.txt",net0.n_0_2_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_5_zneg.txt",net0.n_0_2_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_6_local.txt",net0.n_0_2_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_6_xpos.txt",net0.n_0_2_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_6_xneg.txt",net0.n_0_2_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_6_ypos.txt",net0.n_0_2_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_6_yneg.txt",net0.n_0_2_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_6_zpos.txt",net0.n_0_2_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_6_zneg.txt",net0.n_0_2_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_6_xpos.txt",net0.n_0_2_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_6_xneg.txt",net0.n_0_2_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_6_ypos.txt",net0.n_0_2_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_6_yneg.txt",net0.n_0_2_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_6_zpos.txt",net0.n_0_2_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_6_zneg.txt",net0.n_0_2_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_6_xpos.txt",net0.n_0_2_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_6_xneg.txt",net0.n_0_2_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_6_ypos.txt",net0.n_0_2_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_6_yneg.txt",net0.n_0_2_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_6_zpos.txt",net0.n_0_2_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_6_zneg.txt",net0.n_0_2_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_7_local.txt",net0.n_0_2_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_7_xpos.txt",net0.n_0_2_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_7_xneg.txt",net0.n_0_2_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_7_ypos.txt",net0.n_0_2_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_7_yneg.txt",net0.n_0_2_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_7_zpos.txt",net0.n_0_2_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_2_7_zneg.txt",net0.n_0_2_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_7_xpos.txt",net0.n_0_2_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_7_xneg.txt",net0.n_0_2_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_7_ypos.txt",net0.n_0_2_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_7_yneg.txt",net0.n_0_2_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_7_zpos.txt",net0.n_0_2_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_2_7_zneg.txt",net0.n_0_2_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_7_xpos.txt",net0.n_0_2_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_7_xneg.txt",net0.n_0_2_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_7_ypos.txt",net0.n_0_2_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_7_yneg.txt",net0.n_0_2_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_7_zpos.txt",net0.n_0_2_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_2_7_zneg.txt",net0.n_0_2_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_0_local.txt",net0.n_0_3_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_0_xpos.txt",net0.n_0_3_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_0_xneg.txt",net0.n_0_3_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_0_ypos.txt",net0.n_0_3_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_0_yneg.txt",net0.n_0_3_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_0_zpos.txt",net0.n_0_3_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_0_zneg.txt",net0.n_0_3_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_0_xpos.txt",net0.n_0_3_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_0_xneg.txt",net0.n_0_3_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_0_ypos.txt",net0.n_0_3_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_0_yneg.txt",net0.n_0_3_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_0_zpos.txt",net0.n_0_3_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_0_zneg.txt",net0.n_0_3_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_0_xpos.txt",net0.n_0_3_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_0_xneg.txt",net0.n_0_3_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_0_ypos.txt",net0.n_0_3_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_0_yneg.txt",net0.n_0_3_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_0_zpos.txt",net0.n_0_3_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_0_zneg.txt",net0.n_0_3_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_1_local.txt",net0.n_0_3_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_1_xpos.txt",net0.n_0_3_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_1_xneg.txt",net0.n_0_3_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_1_ypos.txt",net0.n_0_3_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_1_yneg.txt",net0.n_0_3_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_1_zpos.txt",net0.n_0_3_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_1_zneg.txt",net0.n_0_3_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_1_xpos.txt",net0.n_0_3_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_1_xneg.txt",net0.n_0_3_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_1_ypos.txt",net0.n_0_3_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_1_yneg.txt",net0.n_0_3_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_1_zpos.txt",net0.n_0_3_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_1_zneg.txt",net0.n_0_3_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_1_xpos.txt",net0.n_0_3_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_1_xneg.txt",net0.n_0_3_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_1_ypos.txt",net0.n_0_3_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_1_yneg.txt",net0.n_0_3_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_1_zpos.txt",net0.n_0_3_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_1_zneg.txt",net0.n_0_3_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_2_local.txt",net0.n_0_3_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_2_xpos.txt",net0.n_0_3_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_2_xneg.txt",net0.n_0_3_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_2_ypos.txt",net0.n_0_3_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_2_yneg.txt",net0.n_0_3_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_2_zpos.txt",net0.n_0_3_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_2_zneg.txt",net0.n_0_3_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_2_xpos.txt",net0.n_0_3_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_2_xneg.txt",net0.n_0_3_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_2_ypos.txt",net0.n_0_3_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_2_yneg.txt",net0.n_0_3_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_2_zpos.txt",net0.n_0_3_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_2_zneg.txt",net0.n_0_3_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_2_xpos.txt",net0.n_0_3_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_2_xneg.txt",net0.n_0_3_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_2_ypos.txt",net0.n_0_3_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_2_yneg.txt",net0.n_0_3_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_2_zpos.txt",net0.n_0_3_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_2_zneg.txt",net0.n_0_3_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_3_local.txt",net0.n_0_3_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_3_xpos.txt",net0.n_0_3_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_3_xneg.txt",net0.n_0_3_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_3_ypos.txt",net0.n_0_3_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_3_yneg.txt",net0.n_0_3_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_3_zpos.txt",net0.n_0_3_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_3_zneg.txt",net0.n_0_3_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_3_xpos.txt",net0.n_0_3_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_3_xneg.txt",net0.n_0_3_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_3_ypos.txt",net0.n_0_3_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_3_yneg.txt",net0.n_0_3_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_3_zpos.txt",net0.n_0_3_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_3_zneg.txt",net0.n_0_3_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_3_xpos.txt",net0.n_0_3_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_3_xneg.txt",net0.n_0_3_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_3_ypos.txt",net0.n_0_3_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_3_yneg.txt",net0.n_0_3_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_3_zpos.txt",net0.n_0_3_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_3_zneg.txt",net0.n_0_3_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_4_local.txt",net0.n_0_3_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_4_xpos.txt",net0.n_0_3_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_4_xneg.txt",net0.n_0_3_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_4_ypos.txt",net0.n_0_3_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_4_yneg.txt",net0.n_0_3_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_4_zpos.txt",net0.n_0_3_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_4_zneg.txt",net0.n_0_3_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_4_xpos.txt",net0.n_0_3_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_4_xneg.txt",net0.n_0_3_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_4_ypos.txt",net0.n_0_3_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_4_yneg.txt",net0.n_0_3_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_4_zpos.txt",net0.n_0_3_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_4_zneg.txt",net0.n_0_3_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_4_xpos.txt",net0.n_0_3_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_4_xneg.txt",net0.n_0_3_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_4_ypos.txt",net0.n_0_3_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_4_yneg.txt",net0.n_0_3_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_4_zpos.txt",net0.n_0_3_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_4_zneg.txt",net0.n_0_3_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_5_local.txt",net0.n_0_3_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_5_xpos.txt",net0.n_0_3_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_5_xneg.txt",net0.n_0_3_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_5_ypos.txt",net0.n_0_3_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_5_yneg.txt",net0.n_0_3_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_5_zpos.txt",net0.n_0_3_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_5_zneg.txt",net0.n_0_3_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_5_xpos.txt",net0.n_0_3_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_5_xneg.txt",net0.n_0_3_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_5_ypos.txt",net0.n_0_3_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_5_yneg.txt",net0.n_0_3_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_5_zpos.txt",net0.n_0_3_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_5_zneg.txt",net0.n_0_3_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_5_xpos.txt",net0.n_0_3_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_5_xneg.txt",net0.n_0_3_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_5_ypos.txt",net0.n_0_3_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_5_yneg.txt",net0.n_0_3_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_5_zpos.txt",net0.n_0_3_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_5_zneg.txt",net0.n_0_3_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_6_local.txt",net0.n_0_3_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_6_xpos.txt",net0.n_0_3_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_6_xneg.txt",net0.n_0_3_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_6_ypos.txt",net0.n_0_3_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_6_yneg.txt",net0.n_0_3_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_6_zpos.txt",net0.n_0_3_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_6_zneg.txt",net0.n_0_3_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_6_xpos.txt",net0.n_0_3_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_6_xneg.txt",net0.n_0_3_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_6_ypos.txt",net0.n_0_3_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_6_yneg.txt",net0.n_0_3_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_6_zpos.txt",net0.n_0_3_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_6_zneg.txt",net0.n_0_3_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_6_xpos.txt",net0.n_0_3_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_6_xneg.txt",net0.n_0_3_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_6_ypos.txt",net0.n_0_3_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_6_yneg.txt",net0.n_0_3_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_6_zpos.txt",net0.n_0_3_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_6_zneg.txt",net0.n_0_3_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_7_local.txt",net0.n_0_3_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_7_xpos.txt",net0.n_0_3_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_7_xneg.txt",net0.n_0_3_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_7_ypos.txt",net0.n_0_3_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_7_yneg.txt",net0.n_0_3_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_7_zpos.txt",net0.n_0_3_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_3_7_zneg.txt",net0.n_0_3_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_7_xpos.txt",net0.n_0_3_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_7_xneg.txt",net0.n_0_3_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_7_ypos.txt",net0.n_0_3_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_7_yneg.txt",net0.n_0_3_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_7_zpos.txt",net0.n_0_3_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_3_7_zneg.txt",net0.n_0_3_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_7_xpos.txt",net0.n_0_3_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_7_xneg.txt",net0.n_0_3_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_7_ypos.txt",net0.n_0_3_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_7_yneg.txt",net0.n_0_3_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_7_zpos.txt",net0.n_0_3_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_3_7_zneg.txt",net0.n_0_3_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_0_local.txt",net0.n_0_4_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_0_xpos.txt",net0.n_0_4_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_0_xneg.txt",net0.n_0_4_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_0_ypos.txt",net0.n_0_4_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_0_yneg.txt",net0.n_0_4_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_0_zpos.txt",net0.n_0_4_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_0_zneg.txt",net0.n_0_4_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_0_xpos.txt",net0.n_0_4_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_0_xneg.txt",net0.n_0_4_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_0_ypos.txt",net0.n_0_4_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_0_yneg.txt",net0.n_0_4_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_0_zpos.txt",net0.n_0_4_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_0_zneg.txt",net0.n_0_4_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_0_xpos.txt",net0.n_0_4_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_0_xneg.txt",net0.n_0_4_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_0_ypos.txt",net0.n_0_4_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_0_yneg.txt",net0.n_0_4_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_0_zpos.txt",net0.n_0_4_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_0_zneg.txt",net0.n_0_4_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_1_local.txt",net0.n_0_4_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_1_xpos.txt",net0.n_0_4_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_1_xneg.txt",net0.n_0_4_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_1_ypos.txt",net0.n_0_4_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_1_yneg.txt",net0.n_0_4_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_1_zpos.txt",net0.n_0_4_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_1_zneg.txt",net0.n_0_4_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_1_xpos.txt",net0.n_0_4_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_1_xneg.txt",net0.n_0_4_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_1_ypos.txt",net0.n_0_4_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_1_yneg.txt",net0.n_0_4_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_1_zpos.txt",net0.n_0_4_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_1_zneg.txt",net0.n_0_4_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_1_xpos.txt",net0.n_0_4_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_1_xneg.txt",net0.n_0_4_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_1_ypos.txt",net0.n_0_4_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_1_yneg.txt",net0.n_0_4_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_1_zpos.txt",net0.n_0_4_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_1_zneg.txt",net0.n_0_4_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_2_local.txt",net0.n_0_4_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_2_xpos.txt",net0.n_0_4_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_2_xneg.txt",net0.n_0_4_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_2_ypos.txt",net0.n_0_4_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_2_yneg.txt",net0.n_0_4_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_2_zpos.txt",net0.n_0_4_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_2_zneg.txt",net0.n_0_4_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_2_xpos.txt",net0.n_0_4_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_2_xneg.txt",net0.n_0_4_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_2_ypos.txt",net0.n_0_4_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_2_yneg.txt",net0.n_0_4_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_2_zpos.txt",net0.n_0_4_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_2_zneg.txt",net0.n_0_4_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_2_xpos.txt",net0.n_0_4_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_2_xneg.txt",net0.n_0_4_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_2_ypos.txt",net0.n_0_4_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_2_yneg.txt",net0.n_0_4_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_2_zpos.txt",net0.n_0_4_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_2_zneg.txt",net0.n_0_4_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_3_local.txt",net0.n_0_4_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_3_xpos.txt",net0.n_0_4_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_3_xneg.txt",net0.n_0_4_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_3_ypos.txt",net0.n_0_4_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_3_yneg.txt",net0.n_0_4_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_3_zpos.txt",net0.n_0_4_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_3_zneg.txt",net0.n_0_4_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_3_xpos.txt",net0.n_0_4_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_3_xneg.txt",net0.n_0_4_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_3_ypos.txt",net0.n_0_4_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_3_yneg.txt",net0.n_0_4_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_3_zpos.txt",net0.n_0_4_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_3_zneg.txt",net0.n_0_4_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_3_xpos.txt",net0.n_0_4_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_3_xneg.txt",net0.n_0_4_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_3_ypos.txt",net0.n_0_4_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_3_yneg.txt",net0.n_0_4_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_3_zpos.txt",net0.n_0_4_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_3_zneg.txt",net0.n_0_4_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_4_local.txt",net0.n_0_4_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_4_xpos.txt",net0.n_0_4_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_4_xneg.txt",net0.n_0_4_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_4_ypos.txt",net0.n_0_4_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_4_yneg.txt",net0.n_0_4_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_4_zpos.txt",net0.n_0_4_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_4_zneg.txt",net0.n_0_4_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_4_xpos.txt",net0.n_0_4_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_4_xneg.txt",net0.n_0_4_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_4_ypos.txt",net0.n_0_4_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_4_yneg.txt",net0.n_0_4_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_4_zpos.txt",net0.n_0_4_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_4_zneg.txt",net0.n_0_4_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_4_xpos.txt",net0.n_0_4_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_4_xneg.txt",net0.n_0_4_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_4_ypos.txt",net0.n_0_4_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_4_yneg.txt",net0.n_0_4_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_4_zpos.txt",net0.n_0_4_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_4_zneg.txt",net0.n_0_4_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_5_local.txt",net0.n_0_4_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_5_xpos.txt",net0.n_0_4_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_5_xneg.txt",net0.n_0_4_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_5_ypos.txt",net0.n_0_4_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_5_yneg.txt",net0.n_0_4_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_5_zpos.txt",net0.n_0_4_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_5_zneg.txt",net0.n_0_4_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_5_xpos.txt",net0.n_0_4_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_5_xneg.txt",net0.n_0_4_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_5_ypos.txt",net0.n_0_4_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_5_yneg.txt",net0.n_0_4_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_5_zpos.txt",net0.n_0_4_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_5_zneg.txt",net0.n_0_4_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_5_xpos.txt",net0.n_0_4_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_5_xneg.txt",net0.n_0_4_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_5_ypos.txt",net0.n_0_4_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_5_yneg.txt",net0.n_0_4_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_5_zpos.txt",net0.n_0_4_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_5_zneg.txt",net0.n_0_4_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_6_local.txt",net0.n_0_4_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_6_xpos.txt",net0.n_0_4_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_6_xneg.txt",net0.n_0_4_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_6_ypos.txt",net0.n_0_4_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_6_yneg.txt",net0.n_0_4_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_6_zpos.txt",net0.n_0_4_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_6_zneg.txt",net0.n_0_4_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_6_xpos.txt",net0.n_0_4_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_6_xneg.txt",net0.n_0_4_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_6_ypos.txt",net0.n_0_4_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_6_yneg.txt",net0.n_0_4_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_6_zpos.txt",net0.n_0_4_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_6_zneg.txt",net0.n_0_4_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_6_xpos.txt",net0.n_0_4_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_6_xneg.txt",net0.n_0_4_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_6_ypos.txt",net0.n_0_4_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_6_yneg.txt",net0.n_0_4_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_6_zpos.txt",net0.n_0_4_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_6_zneg.txt",net0.n_0_4_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_7_local.txt",net0.n_0_4_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_7_xpos.txt",net0.n_0_4_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_7_xneg.txt",net0.n_0_4_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_7_ypos.txt",net0.n_0_4_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_7_yneg.txt",net0.n_0_4_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_7_zpos.txt",net0.n_0_4_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_4_7_zneg.txt",net0.n_0_4_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_7_xpos.txt",net0.n_0_4_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_7_xneg.txt",net0.n_0_4_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_7_ypos.txt",net0.n_0_4_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_7_yneg.txt",net0.n_0_4_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_7_zpos.txt",net0.n_0_4_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_4_7_zneg.txt",net0.n_0_4_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_7_xpos.txt",net0.n_0_4_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_7_xneg.txt",net0.n_0_4_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_7_ypos.txt",net0.n_0_4_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_7_yneg.txt",net0.n_0_4_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_7_zpos.txt",net0.n_0_4_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_4_7_zneg.txt",net0.n_0_4_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_0_local.txt",net0.n_0_5_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_0_xpos.txt",net0.n_0_5_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_0_xneg.txt",net0.n_0_5_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_0_ypos.txt",net0.n_0_5_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_0_yneg.txt",net0.n_0_5_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_0_zpos.txt",net0.n_0_5_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_0_zneg.txt",net0.n_0_5_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_0_xpos.txt",net0.n_0_5_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_0_xneg.txt",net0.n_0_5_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_0_ypos.txt",net0.n_0_5_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_0_yneg.txt",net0.n_0_5_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_0_zpos.txt",net0.n_0_5_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_0_zneg.txt",net0.n_0_5_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_0_xpos.txt",net0.n_0_5_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_0_xneg.txt",net0.n_0_5_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_0_ypos.txt",net0.n_0_5_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_0_yneg.txt",net0.n_0_5_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_0_zpos.txt",net0.n_0_5_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_0_zneg.txt",net0.n_0_5_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_1_local.txt",net0.n_0_5_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_1_xpos.txt",net0.n_0_5_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_1_xneg.txt",net0.n_0_5_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_1_ypos.txt",net0.n_0_5_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_1_yneg.txt",net0.n_0_5_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_1_zpos.txt",net0.n_0_5_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_1_zneg.txt",net0.n_0_5_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_1_xpos.txt",net0.n_0_5_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_1_xneg.txt",net0.n_0_5_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_1_ypos.txt",net0.n_0_5_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_1_yneg.txt",net0.n_0_5_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_1_zpos.txt",net0.n_0_5_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_1_zneg.txt",net0.n_0_5_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_1_xpos.txt",net0.n_0_5_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_1_xneg.txt",net0.n_0_5_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_1_ypos.txt",net0.n_0_5_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_1_yneg.txt",net0.n_0_5_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_1_zpos.txt",net0.n_0_5_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_1_zneg.txt",net0.n_0_5_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_2_local.txt",net0.n_0_5_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_2_xpos.txt",net0.n_0_5_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_2_xneg.txt",net0.n_0_5_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_2_ypos.txt",net0.n_0_5_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_2_yneg.txt",net0.n_0_5_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_2_zpos.txt",net0.n_0_5_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_2_zneg.txt",net0.n_0_5_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_2_xpos.txt",net0.n_0_5_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_2_xneg.txt",net0.n_0_5_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_2_ypos.txt",net0.n_0_5_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_2_yneg.txt",net0.n_0_5_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_2_zpos.txt",net0.n_0_5_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_2_zneg.txt",net0.n_0_5_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_2_xpos.txt",net0.n_0_5_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_2_xneg.txt",net0.n_0_5_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_2_ypos.txt",net0.n_0_5_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_2_yneg.txt",net0.n_0_5_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_2_zpos.txt",net0.n_0_5_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_2_zneg.txt",net0.n_0_5_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_3_local.txt",net0.n_0_5_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_3_xpos.txt",net0.n_0_5_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_3_xneg.txt",net0.n_0_5_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_3_ypos.txt",net0.n_0_5_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_3_yneg.txt",net0.n_0_5_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_3_zpos.txt",net0.n_0_5_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_3_zneg.txt",net0.n_0_5_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_3_xpos.txt",net0.n_0_5_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_3_xneg.txt",net0.n_0_5_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_3_ypos.txt",net0.n_0_5_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_3_yneg.txt",net0.n_0_5_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_3_zpos.txt",net0.n_0_5_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_3_zneg.txt",net0.n_0_5_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_3_xpos.txt",net0.n_0_5_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_3_xneg.txt",net0.n_0_5_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_3_ypos.txt",net0.n_0_5_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_3_yneg.txt",net0.n_0_5_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_3_zpos.txt",net0.n_0_5_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_3_zneg.txt",net0.n_0_5_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_4_local.txt",net0.n_0_5_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_4_xpos.txt",net0.n_0_5_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_4_xneg.txt",net0.n_0_5_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_4_ypos.txt",net0.n_0_5_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_4_yneg.txt",net0.n_0_5_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_4_zpos.txt",net0.n_0_5_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_4_zneg.txt",net0.n_0_5_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_4_xpos.txt",net0.n_0_5_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_4_xneg.txt",net0.n_0_5_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_4_ypos.txt",net0.n_0_5_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_4_yneg.txt",net0.n_0_5_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_4_zpos.txt",net0.n_0_5_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_4_zneg.txt",net0.n_0_5_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_4_xpos.txt",net0.n_0_5_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_4_xneg.txt",net0.n_0_5_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_4_ypos.txt",net0.n_0_5_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_4_yneg.txt",net0.n_0_5_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_4_zpos.txt",net0.n_0_5_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_4_zneg.txt",net0.n_0_5_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_5_local.txt",net0.n_0_5_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_5_xpos.txt",net0.n_0_5_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_5_xneg.txt",net0.n_0_5_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_5_ypos.txt",net0.n_0_5_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_5_yneg.txt",net0.n_0_5_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_5_zpos.txt",net0.n_0_5_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_5_zneg.txt",net0.n_0_5_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_5_xpos.txt",net0.n_0_5_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_5_xneg.txt",net0.n_0_5_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_5_ypos.txt",net0.n_0_5_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_5_yneg.txt",net0.n_0_5_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_5_zpos.txt",net0.n_0_5_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_5_zneg.txt",net0.n_0_5_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_5_xpos.txt",net0.n_0_5_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_5_xneg.txt",net0.n_0_5_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_5_ypos.txt",net0.n_0_5_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_5_yneg.txt",net0.n_0_5_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_5_zpos.txt",net0.n_0_5_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_5_zneg.txt",net0.n_0_5_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_6_local.txt",net0.n_0_5_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_6_xpos.txt",net0.n_0_5_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_6_xneg.txt",net0.n_0_5_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_6_ypos.txt",net0.n_0_5_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_6_yneg.txt",net0.n_0_5_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_6_zpos.txt",net0.n_0_5_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_6_zneg.txt",net0.n_0_5_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_6_xpos.txt",net0.n_0_5_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_6_xneg.txt",net0.n_0_5_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_6_ypos.txt",net0.n_0_5_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_6_yneg.txt",net0.n_0_5_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_6_zpos.txt",net0.n_0_5_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_6_zneg.txt",net0.n_0_5_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_6_xpos.txt",net0.n_0_5_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_6_xneg.txt",net0.n_0_5_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_6_ypos.txt",net0.n_0_5_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_6_yneg.txt",net0.n_0_5_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_6_zpos.txt",net0.n_0_5_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_6_zneg.txt",net0.n_0_5_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_7_local.txt",net0.n_0_5_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_7_xpos.txt",net0.n_0_5_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_7_xneg.txt",net0.n_0_5_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_7_ypos.txt",net0.n_0_5_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_7_yneg.txt",net0.n_0_5_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_7_zpos.txt",net0.n_0_5_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_5_7_zneg.txt",net0.n_0_5_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_7_xpos.txt",net0.n_0_5_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_7_xneg.txt",net0.n_0_5_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_7_ypos.txt",net0.n_0_5_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_7_yneg.txt",net0.n_0_5_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_7_zpos.txt",net0.n_0_5_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_5_7_zneg.txt",net0.n_0_5_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_7_xpos.txt",net0.n_0_5_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_7_xneg.txt",net0.n_0_5_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_7_ypos.txt",net0.n_0_5_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_7_yneg.txt",net0.n_0_5_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_7_zpos.txt",net0.n_0_5_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_5_7_zneg.txt",net0.n_0_5_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_0_local.txt",net0.n_0_6_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_0_xpos.txt",net0.n_0_6_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_0_xneg.txt",net0.n_0_6_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_0_ypos.txt",net0.n_0_6_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_0_yneg.txt",net0.n_0_6_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_0_zpos.txt",net0.n_0_6_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_0_zneg.txt",net0.n_0_6_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_0_xpos.txt",net0.n_0_6_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_0_xneg.txt",net0.n_0_6_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_0_ypos.txt",net0.n_0_6_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_0_yneg.txt",net0.n_0_6_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_0_zpos.txt",net0.n_0_6_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_0_zneg.txt",net0.n_0_6_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_0_xpos.txt",net0.n_0_6_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_0_xneg.txt",net0.n_0_6_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_0_ypos.txt",net0.n_0_6_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_0_yneg.txt",net0.n_0_6_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_0_zpos.txt",net0.n_0_6_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_0_zneg.txt",net0.n_0_6_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_1_local.txt",net0.n_0_6_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_1_xpos.txt",net0.n_0_6_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_1_xneg.txt",net0.n_0_6_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_1_ypos.txt",net0.n_0_6_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_1_yneg.txt",net0.n_0_6_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_1_zpos.txt",net0.n_0_6_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_1_zneg.txt",net0.n_0_6_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_1_xpos.txt",net0.n_0_6_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_1_xneg.txt",net0.n_0_6_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_1_ypos.txt",net0.n_0_6_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_1_yneg.txt",net0.n_0_6_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_1_zpos.txt",net0.n_0_6_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_1_zneg.txt",net0.n_0_6_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_1_xpos.txt",net0.n_0_6_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_1_xneg.txt",net0.n_0_6_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_1_ypos.txt",net0.n_0_6_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_1_yneg.txt",net0.n_0_6_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_1_zpos.txt",net0.n_0_6_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_1_zneg.txt",net0.n_0_6_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_2_local.txt",net0.n_0_6_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_2_xpos.txt",net0.n_0_6_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_2_xneg.txt",net0.n_0_6_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_2_ypos.txt",net0.n_0_6_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_2_yneg.txt",net0.n_0_6_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_2_zpos.txt",net0.n_0_6_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_2_zneg.txt",net0.n_0_6_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_2_xpos.txt",net0.n_0_6_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_2_xneg.txt",net0.n_0_6_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_2_ypos.txt",net0.n_0_6_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_2_yneg.txt",net0.n_0_6_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_2_zpos.txt",net0.n_0_6_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_2_zneg.txt",net0.n_0_6_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_2_xpos.txt",net0.n_0_6_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_2_xneg.txt",net0.n_0_6_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_2_ypos.txt",net0.n_0_6_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_2_yneg.txt",net0.n_0_6_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_2_zpos.txt",net0.n_0_6_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_2_zneg.txt",net0.n_0_6_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_3_local.txt",net0.n_0_6_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_3_xpos.txt",net0.n_0_6_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_3_xneg.txt",net0.n_0_6_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_3_ypos.txt",net0.n_0_6_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_3_yneg.txt",net0.n_0_6_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_3_zpos.txt",net0.n_0_6_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_3_zneg.txt",net0.n_0_6_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_3_xpos.txt",net0.n_0_6_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_3_xneg.txt",net0.n_0_6_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_3_ypos.txt",net0.n_0_6_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_3_yneg.txt",net0.n_0_6_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_3_zpos.txt",net0.n_0_6_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_3_zneg.txt",net0.n_0_6_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_3_xpos.txt",net0.n_0_6_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_3_xneg.txt",net0.n_0_6_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_3_ypos.txt",net0.n_0_6_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_3_yneg.txt",net0.n_0_6_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_3_zpos.txt",net0.n_0_6_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_3_zneg.txt",net0.n_0_6_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_4_local.txt",net0.n_0_6_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_4_xpos.txt",net0.n_0_6_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_4_xneg.txt",net0.n_0_6_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_4_ypos.txt",net0.n_0_6_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_4_yneg.txt",net0.n_0_6_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_4_zpos.txt",net0.n_0_6_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_4_zneg.txt",net0.n_0_6_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_4_xpos.txt",net0.n_0_6_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_4_xneg.txt",net0.n_0_6_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_4_ypos.txt",net0.n_0_6_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_4_yneg.txt",net0.n_0_6_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_4_zpos.txt",net0.n_0_6_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_4_zneg.txt",net0.n_0_6_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_4_xpos.txt",net0.n_0_6_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_4_xneg.txt",net0.n_0_6_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_4_ypos.txt",net0.n_0_6_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_4_yneg.txt",net0.n_0_6_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_4_zpos.txt",net0.n_0_6_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_4_zneg.txt",net0.n_0_6_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_5_local.txt",net0.n_0_6_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_5_xpos.txt",net0.n_0_6_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_5_xneg.txt",net0.n_0_6_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_5_ypos.txt",net0.n_0_6_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_5_yneg.txt",net0.n_0_6_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_5_zpos.txt",net0.n_0_6_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_5_zneg.txt",net0.n_0_6_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_5_xpos.txt",net0.n_0_6_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_5_xneg.txt",net0.n_0_6_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_5_ypos.txt",net0.n_0_6_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_5_yneg.txt",net0.n_0_6_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_5_zpos.txt",net0.n_0_6_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_5_zneg.txt",net0.n_0_6_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_5_xpos.txt",net0.n_0_6_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_5_xneg.txt",net0.n_0_6_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_5_ypos.txt",net0.n_0_6_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_5_yneg.txt",net0.n_0_6_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_5_zpos.txt",net0.n_0_6_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_5_zneg.txt",net0.n_0_6_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_6_local.txt",net0.n_0_6_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_6_xpos.txt",net0.n_0_6_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_6_xneg.txt",net0.n_0_6_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_6_ypos.txt",net0.n_0_6_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_6_yneg.txt",net0.n_0_6_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_6_zpos.txt",net0.n_0_6_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_6_zneg.txt",net0.n_0_6_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_6_xpos.txt",net0.n_0_6_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_6_xneg.txt",net0.n_0_6_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_6_ypos.txt",net0.n_0_6_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_6_yneg.txt",net0.n_0_6_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_6_zpos.txt",net0.n_0_6_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_6_zneg.txt",net0.n_0_6_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_6_xpos.txt",net0.n_0_6_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_6_xneg.txt",net0.n_0_6_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_6_ypos.txt",net0.n_0_6_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_6_yneg.txt",net0.n_0_6_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_6_zpos.txt",net0.n_0_6_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_6_zneg.txt",net0.n_0_6_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_7_local.txt",net0.n_0_6_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_7_xpos.txt",net0.n_0_6_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_7_xneg.txt",net0.n_0_6_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_7_ypos.txt",net0.n_0_6_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_7_yneg.txt",net0.n_0_6_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_7_zpos.txt",net0.n_0_6_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_6_7_zneg.txt",net0.n_0_6_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_7_xpos.txt",net0.n_0_6_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_7_xneg.txt",net0.n_0_6_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_7_ypos.txt",net0.n_0_6_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_7_yneg.txt",net0.n_0_6_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_7_zpos.txt",net0.n_0_6_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_6_7_zneg.txt",net0.n_0_6_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_7_xpos.txt",net0.n_0_6_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_7_xneg.txt",net0.n_0_6_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_7_ypos.txt",net0.n_0_6_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_7_yneg.txt",net0.n_0_6_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_7_zpos.txt",net0.n_0_6_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_6_7_zneg.txt",net0.n_0_6_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_0_local.txt",net0.n_0_7_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_0_xpos.txt",net0.n_0_7_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_0_xneg.txt",net0.n_0_7_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_0_ypos.txt",net0.n_0_7_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_0_yneg.txt",net0.n_0_7_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_0_zpos.txt",net0.n_0_7_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_0_zneg.txt",net0.n_0_7_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_0_xpos.txt",net0.n_0_7_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_0_xneg.txt",net0.n_0_7_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_0_ypos.txt",net0.n_0_7_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_0_yneg.txt",net0.n_0_7_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_0_zpos.txt",net0.n_0_7_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_0_zneg.txt",net0.n_0_7_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_0_xpos.txt",net0.n_0_7_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_0_xneg.txt",net0.n_0_7_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_0_ypos.txt",net0.n_0_7_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_0_yneg.txt",net0.n_0_7_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_0_zpos.txt",net0.n_0_7_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_0_zneg.txt",net0.n_0_7_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_1_local.txt",net0.n_0_7_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_1_xpos.txt",net0.n_0_7_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_1_xneg.txt",net0.n_0_7_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_1_ypos.txt",net0.n_0_7_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_1_yneg.txt",net0.n_0_7_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_1_zpos.txt",net0.n_0_7_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_1_zneg.txt",net0.n_0_7_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_1_xpos.txt",net0.n_0_7_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_1_xneg.txt",net0.n_0_7_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_1_ypos.txt",net0.n_0_7_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_1_yneg.txt",net0.n_0_7_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_1_zpos.txt",net0.n_0_7_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_1_zneg.txt",net0.n_0_7_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_1_xpos.txt",net0.n_0_7_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_1_xneg.txt",net0.n_0_7_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_1_ypos.txt",net0.n_0_7_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_1_yneg.txt",net0.n_0_7_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_1_zpos.txt",net0.n_0_7_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_1_zneg.txt",net0.n_0_7_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_2_local.txt",net0.n_0_7_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_2_xpos.txt",net0.n_0_7_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_2_xneg.txt",net0.n_0_7_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_2_ypos.txt",net0.n_0_7_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_2_yneg.txt",net0.n_0_7_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_2_zpos.txt",net0.n_0_7_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_2_zneg.txt",net0.n_0_7_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_2_xpos.txt",net0.n_0_7_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_2_xneg.txt",net0.n_0_7_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_2_ypos.txt",net0.n_0_7_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_2_yneg.txt",net0.n_0_7_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_2_zpos.txt",net0.n_0_7_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_2_zneg.txt",net0.n_0_7_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_2_xpos.txt",net0.n_0_7_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_2_xneg.txt",net0.n_0_7_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_2_ypos.txt",net0.n_0_7_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_2_yneg.txt",net0.n_0_7_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_2_zpos.txt",net0.n_0_7_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_2_zneg.txt",net0.n_0_7_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_3_local.txt",net0.n_0_7_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_3_xpos.txt",net0.n_0_7_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_3_xneg.txt",net0.n_0_7_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_3_ypos.txt",net0.n_0_7_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_3_yneg.txt",net0.n_0_7_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_3_zpos.txt",net0.n_0_7_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_3_zneg.txt",net0.n_0_7_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_3_xpos.txt",net0.n_0_7_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_3_xneg.txt",net0.n_0_7_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_3_ypos.txt",net0.n_0_7_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_3_yneg.txt",net0.n_0_7_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_3_zpos.txt",net0.n_0_7_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_3_zneg.txt",net0.n_0_7_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_3_xpos.txt",net0.n_0_7_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_3_xneg.txt",net0.n_0_7_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_3_ypos.txt",net0.n_0_7_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_3_yneg.txt",net0.n_0_7_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_3_zpos.txt",net0.n_0_7_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_3_zneg.txt",net0.n_0_7_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_4_local.txt",net0.n_0_7_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_4_xpos.txt",net0.n_0_7_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_4_xneg.txt",net0.n_0_7_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_4_ypos.txt",net0.n_0_7_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_4_yneg.txt",net0.n_0_7_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_4_zpos.txt",net0.n_0_7_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_4_zneg.txt",net0.n_0_7_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_4_xpos.txt",net0.n_0_7_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_4_xneg.txt",net0.n_0_7_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_4_ypos.txt",net0.n_0_7_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_4_yneg.txt",net0.n_0_7_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_4_zpos.txt",net0.n_0_7_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_4_zneg.txt",net0.n_0_7_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_4_xpos.txt",net0.n_0_7_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_4_xneg.txt",net0.n_0_7_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_4_ypos.txt",net0.n_0_7_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_4_yneg.txt",net0.n_0_7_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_4_zpos.txt",net0.n_0_7_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_4_zneg.txt",net0.n_0_7_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_5_local.txt",net0.n_0_7_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_5_xpos.txt",net0.n_0_7_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_5_xneg.txt",net0.n_0_7_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_5_ypos.txt",net0.n_0_7_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_5_yneg.txt",net0.n_0_7_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_5_zpos.txt",net0.n_0_7_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_5_zneg.txt",net0.n_0_7_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_5_xpos.txt",net0.n_0_7_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_5_xneg.txt",net0.n_0_7_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_5_ypos.txt",net0.n_0_7_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_5_yneg.txt",net0.n_0_7_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_5_zpos.txt",net0.n_0_7_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_5_zneg.txt",net0.n_0_7_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_5_xpos.txt",net0.n_0_7_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_5_xneg.txt",net0.n_0_7_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_5_ypos.txt",net0.n_0_7_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_5_yneg.txt",net0.n_0_7_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_5_zpos.txt",net0.n_0_7_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_5_zneg.txt",net0.n_0_7_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_6_local.txt",net0.n_0_7_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_6_xpos.txt",net0.n_0_7_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_6_xneg.txt",net0.n_0_7_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_6_ypos.txt",net0.n_0_7_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_6_yneg.txt",net0.n_0_7_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_6_zpos.txt",net0.n_0_7_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_6_zneg.txt",net0.n_0_7_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_6_xpos.txt",net0.n_0_7_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_6_xneg.txt",net0.n_0_7_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_6_ypos.txt",net0.n_0_7_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_6_yneg.txt",net0.n_0_7_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_6_zpos.txt",net0.n_0_7_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_6_zneg.txt",net0.n_0_7_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_6_xpos.txt",net0.n_0_7_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_6_xneg.txt",net0.n_0_7_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_6_ypos.txt",net0.n_0_7_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_6_yneg.txt",net0.n_0_7_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_6_zpos.txt",net0.n_0_7_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_6_zneg.txt",net0.n_0_7_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_7_local.txt",net0.n_0_7_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_7_xpos.txt",net0.n_0_7_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_7_xneg.txt",net0.n_0_7_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_7_ypos.txt",net0.n_0_7_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_7_yneg.txt",net0.n_0_7_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_7_zpos.txt",net0.n_0_7_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_0_7_7_zneg.txt",net0.n_0_7_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_7_xpos.txt",net0.n_0_7_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_7_xneg.txt",net0.n_0_7_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_7_ypos.txt",net0.n_0_7_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_7_yneg.txt",net0.n_0_7_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_7_zpos.txt",net0.n_0_7_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_0_7_7_zneg.txt",net0.n_0_7_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_7_xpos.txt",net0.n_0_7_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_7_xneg.txt",net0.n_0_7_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_7_ypos.txt",net0.n_0_7_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_7_yneg.txt",net0.n_0_7_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_7_zpos.txt",net0.n_0_7_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_0_7_7_zneg.txt",net0.n_0_7_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_0_local.txt",net0.n_1_0_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_0_xpos.txt",net0.n_1_0_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_0_xneg.txt",net0.n_1_0_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_0_ypos.txt",net0.n_1_0_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_0_yneg.txt",net0.n_1_0_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_0_zpos.txt",net0.n_1_0_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_0_zneg.txt",net0.n_1_0_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_0_xpos.txt",net0.n_1_0_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_0_xneg.txt",net0.n_1_0_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_0_ypos.txt",net0.n_1_0_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_0_yneg.txt",net0.n_1_0_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_0_zpos.txt",net0.n_1_0_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_0_zneg.txt",net0.n_1_0_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_0_xpos.txt",net0.n_1_0_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_0_xneg.txt",net0.n_1_0_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_0_ypos.txt",net0.n_1_0_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_0_yneg.txt",net0.n_1_0_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_0_zpos.txt",net0.n_1_0_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_0_zneg.txt",net0.n_1_0_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_1_local.txt",net0.n_1_0_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_1_xpos.txt",net0.n_1_0_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_1_xneg.txt",net0.n_1_0_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_1_ypos.txt",net0.n_1_0_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_1_yneg.txt",net0.n_1_0_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_1_zpos.txt",net0.n_1_0_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_1_zneg.txt",net0.n_1_0_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_1_xpos.txt",net0.n_1_0_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_1_xneg.txt",net0.n_1_0_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_1_ypos.txt",net0.n_1_0_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_1_yneg.txt",net0.n_1_0_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_1_zpos.txt",net0.n_1_0_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_1_zneg.txt",net0.n_1_0_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_1_xpos.txt",net0.n_1_0_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_1_xneg.txt",net0.n_1_0_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_1_ypos.txt",net0.n_1_0_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_1_yneg.txt",net0.n_1_0_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_1_zpos.txt",net0.n_1_0_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_1_zneg.txt",net0.n_1_0_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_2_local.txt",net0.n_1_0_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_2_xpos.txt",net0.n_1_0_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_2_xneg.txt",net0.n_1_0_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_2_ypos.txt",net0.n_1_0_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_2_yneg.txt",net0.n_1_0_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_2_zpos.txt",net0.n_1_0_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_2_zneg.txt",net0.n_1_0_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_2_xpos.txt",net0.n_1_0_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_2_xneg.txt",net0.n_1_0_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_2_ypos.txt",net0.n_1_0_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_2_yneg.txt",net0.n_1_0_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_2_zpos.txt",net0.n_1_0_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_2_zneg.txt",net0.n_1_0_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_2_xpos.txt",net0.n_1_0_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_2_xneg.txt",net0.n_1_0_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_2_ypos.txt",net0.n_1_0_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_2_yneg.txt",net0.n_1_0_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_2_zpos.txt",net0.n_1_0_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_2_zneg.txt",net0.n_1_0_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_3_local.txt",net0.n_1_0_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_3_xpos.txt",net0.n_1_0_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_3_xneg.txt",net0.n_1_0_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_3_ypos.txt",net0.n_1_0_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_3_yneg.txt",net0.n_1_0_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_3_zpos.txt",net0.n_1_0_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_3_zneg.txt",net0.n_1_0_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_3_xpos.txt",net0.n_1_0_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_3_xneg.txt",net0.n_1_0_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_3_ypos.txt",net0.n_1_0_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_3_yneg.txt",net0.n_1_0_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_3_zpos.txt",net0.n_1_0_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_3_zneg.txt",net0.n_1_0_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_3_xpos.txt",net0.n_1_0_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_3_xneg.txt",net0.n_1_0_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_3_ypos.txt",net0.n_1_0_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_3_yneg.txt",net0.n_1_0_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_3_zpos.txt",net0.n_1_0_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_3_zneg.txt",net0.n_1_0_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_4_local.txt",net0.n_1_0_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_4_xpos.txt",net0.n_1_0_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_4_xneg.txt",net0.n_1_0_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_4_ypos.txt",net0.n_1_0_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_4_yneg.txt",net0.n_1_0_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_4_zpos.txt",net0.n_1_0_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_4_zneg.txt",net0.n_1_0_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_4_xpos.txt",net0.n_1_0_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_4_xneg.txt",net0.n_1_0_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_4_ypos.txt",net0.n_1_0_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_4_yneg.txt",net0.n_1_0_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_4_zpos.txt",net0.n_1_0_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_4_zneg.txt",net0.n_1_0_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_4_xpos.txt",net0.n_1_0_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_4_xneg.txt",net0.n_1_0_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_4_ypos.txt",net0.n_1_0_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_4_yneg.txt",net0.n_1_0_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_4_zpos.txt",net0.n_1_0_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_4_zneg.txt",net0.n_1_0_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_5_local.txt",net0.n_1_0_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_5_xpos.txt",net0.n_1_0_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_5_xneg.txt",net0.n_1_0_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_5_ypos.txt",net0.n_1_0_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_5_yneg.txt",net0.n_1_0_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_5_zpos.txt",net0.n_1_0_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_5_zneg.txt",net0.n_1_0_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_5_xpos.txt",net0.n_1_0_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_5_xneg.txt",net0.n_1_0_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_5_ypos.txt",net0.n_1_0_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_5_yneg.txt",net0.n_1_0_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_5_zpos.txt",net0.n_1_0_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_5_zneg.txt",net0.n_1_0_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_5_xpos.txt",net0.n_1_0_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_5_xneg.txt",net0.n_1_0_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_5_ypos.txt",net0.n_1_0_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_5_yneg.txt",net0.n_1_0_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_5_zpos.txt",net0.n_1_0_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_5_zneg.txt",net0.n_1_0_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_6_local.txt",net0.n_1_0_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_6_xpos.txt",net0.n_1_0_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_6_xneg.txt",net0.n_1_0_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_6_ypos.txt",net0.n_1_0_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_6_yneg.txt",net0.n_1_0_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_6_zpos.txt",net0.n_1_0_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_6_zneg.txt",net0.n_1_0_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_6_xpos.txt",net0.n_1_0_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_6_xneg.txt",net0.n_1_0_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_6_ypos.txt",net0.n_1_0_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_6_yneg.txt",net0.n_1_0_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_6_zpos.txt",net0.n_1_0_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_6_zneg.txt",net0.n_1_0_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_6_xpos.txt",net0.n_1_0_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_6_xneg.txt",net0.n_1_0_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_6_ypos.txt",net0.n_1_0_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_6_yneg.txt",net0.n_1_0_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_6_zpos.txt",net0.n_1_0_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_6_zneg.txt",net0.n_1_0_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_7_local.txt",net0.n_1_0_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_7_xpos.txt",net0.n_1_0_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_7_xneg.txt",net0.n_1_0_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_7_ypos.txt",net0.n_1_0_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_7_yneg.txt",net0.n_1_0_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_7_zpos.txt",net0.n_1_0_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_0_7_zneg.txt",net0.n_1_0_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_7_xpos.txt",net0.n_1_0_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_7_xneg.txt",net0.n_1_0_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_7_ypos.txt",net0.n_1_0_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_7_yneg.txt",net0.n_1_0_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_7_zpos.txt",net0.n_1_0_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_0_7_zneg.txt",net0.n_1_0_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_7_xpos.txt",net0.n_1_0_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_7_xneg.txt",net0.n_1_0_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_7_ypos.txt",net0.n_1_0_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_7_yneg.txt",net0.n_1_0_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_7_zpos.txt",net0.n_1_0_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_0_7_zneg.txt",net0.n_1_0_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_0_local.txt",net0.n_1_1_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_0_xpos.txt",net0.n_1_1_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_0_xneg.txt",net0.n_1_1_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_0_ypos.txt",net0.n_1_1_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_0_yneg.txt",net0.n_1_1_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_0_zpos.txt",net0.n_1_1_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_0_zneg.txt",net0.n_1_1_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_0_xpos.txt",net0.n_1_1_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_0_xneg.txt",net0.n_1_1_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_0_ypos.txt",net0.n_1_1_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_0_yneg.txt",net0.n_1_1_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_0_zpos.txt",net0.n_1_1_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_0_zneg.txt",net0.n_1_1_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_0_xpos.txt",net0.n_1_1_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_0_xneg.txt",net0.n_1_1_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_0_ypos.txt",net0.n_1_1_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_0_yneg.txt",net0.n_1_1_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_0_zpos.txt",net0.n_1_1_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_0_zneg.txt",net0.n_1_1_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_1_local.txt",net0.n_1_1_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_1_xpos.txt",net0.n_1_1_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_1_xneg.txt",net0.n_1_1_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_1_ypos.txt",net0.n_1_1_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_1_yneg.txt",net0.n_1_1_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_1_zpos.txt",net0.n_1_1_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_1_zneg.txt",net0.n_1_1_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_1_xpos.txt",net0.n_1_1_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_1_xneg.txt",net0.n_1_1_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_1_ypos.txt",net0.n_1_1_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_1_yneg.txt",net0.n_1_1_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_1_zpos.txt",net0.n_1_1_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_1_zneg.txt",net0.n_1_1_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_1_xpos.txt",net0.n_1_1_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_1_xneg.txt",net0.n_1_1_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_1_ypos.txt",net0.n_1_1_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_1_yneg.txt",net0.n_1_1_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_1_zpos.txt",net0.n_1_1_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_1_zneg.txt",net0.n_1_1_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_2_local.txt",net0.n_1_1_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_2_xpos.txt",net0.n_1_1_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_2_xneg.txt",net0.n_1_1_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_2_ypos.txt",net0.n_1_1_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_2_yneg.txt",net0.n_1_1_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_2_zpos.txt",net0.n_1_1_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_2_zneg.txt",net0.n_1_1_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_2_xpos.txt",net0.n_1_1_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_2_xneg.txt",net0.n_1_1_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_2_ypos.txt",net0.n_1_1_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_2_yneg.txt",net0.n_1_1_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_2_zpos.txt",net0.n_1_1_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_2_zneg.txt",net0.n_1_1_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_2_xpos.txt",net0.n_1_1_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_2_xneg.txt",net0.n_1_1_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_2_ypos.txt",net0.n_1_1_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_2_yneg.txt",net0.n_1_1_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_2_zpos.txt",net0.n_1_1_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_2_zneg.txt",net0.n_1_1_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_3_local.txt",net0.n_1_1_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_3_xpos.txt",net0.n_1_1_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_3_xneg.txt",net0.n_1_1_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_3_ypos.txt",net0.n_1_1_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_3_yneg.txt",net0.n_1_1_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_3_zpos.txt",net0.n_1_1_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_3_zneg.txt",net0.n_1_1_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_3_xpos.txt",net0.n_1_1_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_3_xneg.txt",net0.n_1_1_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_3_ypos.txt",net0.n_1_1_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_3_yneg.txt",net0.n_1_1_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_3_zpos.txt",net0.n_1_1_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_3_zneg.txt",net0.n_1_1_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_3_xpos.txt",net0.n_1_1_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_3_xneg.txt",net0.n_1_1_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_3_ypos.txt",net0.n_1_1_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_3_yneg.txt",net0.n_1_1_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_3_zpos.txt",net0.n_1_1_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_3_zneg.txt",net0.n_1_1_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_4_local.txt",net0.n_1_1_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_4_xpos.txt",net0.n_1_1_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_4_xneg.txt",net0.n_1_1_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_4_ypos.txt",net0.n_1_1_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_4_yneg.txt",net0.n_1_1_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_4_zpos.txt",net0.n_1_1_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_4_zneg.txt",net0.n_1_1_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_4_xpos.txt",net0.n_1_1_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_4_xneg.txt",net0.n_1_1_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_4_ypos.txt",net0.n_1_1_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_4_yneg.txt",net0.n_1_1_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_4_zpos.txt",net0.n_1_1_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_4_zneg.txt",net0.n_1_1_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_4_xpos.txt",net0.n_1_1_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_4_xneg.txt",net0.n_1_1_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_4_ypos.txt",net0.n_1_1_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_4_yneg.txt",net0.n_1_1_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_4_zpos.txt",net0.n_1_1_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_4_zneg.txt",net0.n_1_1_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_5_local.txt",net0.n_1_1_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_5_xpos.txt",net0.n_1_1_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_5_xneg.txt",net0.n_1_1_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_5_ypos.txt",net0.n_1_1_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_5_yneg.txt",net0.n_1_1_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_5_zpos.txt",net0.n_1_1_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_5_zneg.txt",net0.n_1_1_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_5_xpos.txt",net0.n_1_1_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_5_xneg.txt",net0.n_1_1_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_5_ypos.txt",net0.n_1_1_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_5_yneg.txt",net0.n_1_1_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_5_zpos.txt",net0.n_1_1_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_5_zneg.txt",net0.n_1_1_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_5_xpos.txt",net0.n_1_1_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_5_xneg.txt",net0.n_1_1_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_5_ypos.txt",net0.n_1_1_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_5_yneg.txt",net0.n_1_1_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_5_zpos.txt",net0.n_1_1_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_5_zneg.txt",net0.n_1_1_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_6_local.txt",net0.n_1_1_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_6_xpos.txt",net0.n_1_1_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_6_xneg.txt",net0.n_1_1_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_6_ypos.txt",net0.n_1_1_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_6_yneg.txt",net0.n_1_1_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_6_zpos.txt",net0.n_1_1_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_6_zneg.txt",net0.n_1_1_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_6_xpos.txt",net0.n_1_1_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_6_xneg.txt",net0.n_1_1_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_6_ypos.txt",net0.n_1_1_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_6_yneg.txt",net0.n_1_1_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_6_zpos.txt",net0.n_1_1_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_6_zneg.txt",net0.n_1_1_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_6_xpos.txt",net0.n_1_1_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_6_xneg.txt",net0.n_1_1_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_6_ypos.txt",net0.n_1_1_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_6_yneg.txt",net0.n_1_1_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_6_zpos.txt",net0.n_1_1_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_6_zneg.txt",net0.n_1_1_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_7_local.txt",net0.n_1_1_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_7_xpos.txt",net0.n_1_1_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_7_xneg.txt",net0.n_1_1_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_7_ypos.txt",net0.n_1_1_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_7_yneg.txt",net0.n_1_1_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_7_zpos.txt",net0.n_1_1_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_1_7_zneg.txt",net0.n_1_1_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_7_xpos.txt",net0.n_1_1_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_7_xneg.txt",net0.n_1_1_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_7_ypos.txt",net0.n_1_1_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_7_yneg.txt",net0.n_1_1_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_7_zpos.txt",net0.n_1_1_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_1_7_zneg.txt",net0.n_1_1_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_7_xpos.txt",net0.n_1_1_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_7_xneg.txt",net0.n_1_1_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_7_ypos.txt",net0.n_1_1_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_7_yneg.txt",net0.n_1_1_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_7_zpos.txt",net0.n_1_1_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_1_7_zneg.txt",net0.n_1_1_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_0_local.txt",net0.n_1_2_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_0_xpos.txt",net0.n_1_2_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_0_xneg.txt",net0.n_1_2_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_0_ypos.txt",net0.n_1_2_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_0_yneg.txt",net0.n_1_2_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_0_zpos.txt",net0.n_1_2_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_0_zneg.txt",net0.n_1_2_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_0_xpos.txt",net0.n_1_2_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_0_xneg.txt",net0.n_1_2_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_0_ypos.txt",net0.n_1_2_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_0_yneg.txt",net0.n_1_2_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_0_zpos.txt",net0.n_1_2_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_0_zneg.txt",net0.n_1_2_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_0_xpos.txt",net0.n_1_2_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_0_xneg.txt",net0.n_1_2_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_0_ypos.txt",net0.n_1_2_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_0_yneg.txt",net0.n_1_2_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_0_zpos.txt",net0.n_1_2_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_0_zneg.txt",net0.n_1_2_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_1_local.txt",net0.n_1_2_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_1_xpos.txt",net0.n_1_2_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_1_xneg.txt",net0.n_1_2_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_1_ypos.txt",net0.n_1_2_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_1_yneg.txt",net0.n_1_2_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_1_zpos.txt",net0.n_1_2_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_1_zneg.txt",net0.n_1_2_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_1_xpos.txt",net0.n_1_2_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_1_xneg.txt",net0.n_1_2_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_1_ypos.txt",net0.n_1_2_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_1_yneg.txt",net0.n_1_2_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_1_zpos.txt",net0.n_1_2_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_1_zneg.txt",net0.n_1_2_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_1_xpos.txt",net0.n_1_2_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_1_xneg.txt",net0.n_1_2_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_1_ypos.txt",net0.n_1_2_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_1_yneg.txt",net0.n_1_2_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_1_zpos.txt",net0.n_1_2_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_1_zneg.txt",net0.n_1_2_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_2_local.txt",net0.n_1_2_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_2_xpos.txt",net0.n_1_2_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_2_xneg.txt",net0.n_1_2_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_2_ypos.txt",net0.n_1_2_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_2_yneg.txt",net0.n_1_2_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_2_zpos.txt",net0.n_1_2_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_2_zneg.txt",net0.n_1_2_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_2_xpos.txt",net0.n_1_2_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_2_xneg.txt",net0.n_1_2_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_2_ypos.txt",net0.n_1_2_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_2_yneg.txt",net0.n_1_2_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_2_zpos.txt",net0.n_1_2_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_2_zneg.txt",net0.n_1_2_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_2_xpos.txt",net0.n_1_2_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_2_xneg.txt",net0.n_1_2_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_2_ypos.txt",net0.n_1_2_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_2_yneg.txt",net0.n_1_2_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_2_zpos.txt",net0.n_1_2_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_2_zneg.txt",net0.n_1_2_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_3_local.txt",net0.n_1_2_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_3_xpos.txt",net0.n_1_2_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_3_xneg.txt",net0.n_1_2_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_3_ypos.txt",net0.n_1_2_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_3_yneg.txt",net0.n_1_2_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_3_zpos.txt",net0.n_1_2_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_3_zneg.txt",net0.n_1_2_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_3_xpos.txt",net0.n_1_2_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_3_xneg.txt",net0.n_1_2_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_3_ypos.txt",net0.n_1_2_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_3_yneg.txt",net0.n_1_2_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_3_zpos.txt",net0.n_1_2_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_3_zneg.txt",net0.n_1_2_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_3_xpos.txt",net0.n_1_2_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_3_xneg.txt",net0.n_1_2_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_3_ypos.txt",net0.n_1_2_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_3_yneg.txt",net0.n_1_2_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_3_zpos.txt",net0.n_1_2_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_3_zneg.txt",net0.n_1_2_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_4_local.txt",net0.n_1_2_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_4_xpos.txt",net0.n_1_2_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_4_xneg.txt",net0.n_1_2_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_4_ypos.txt",net0.n_1_2_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_4_yneg.txt",net0.n_1_2_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_4_zpos.txt",net0.n_1_2_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_4_zneg.txt",net0.n_1_2_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_4_xpos.txt",net0.n_1_2_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_4_xneg.txt",net0.n_1_2_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_4_ypos.txt",net0.n_1_2_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_4_yneg.txt",net0.n_1_2_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_4_zpos.txt",net0.n_1_2_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_4_zneg.txt",net0.n_1_2_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_4_xpos.txt",net0.n_1_2_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_4_xneg.txt",net0.n_1_2_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_4_ypos.txt",net0.n_1_2_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_4_yneg.txt",net0.n_1_2_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_4_zpos.txt",net0.n_1_2_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_4_zneg.txt",net0.n_1_2_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_5_local.txt",net0.n_1_2_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_5_xpos.txt",net0.n_1_2_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_5_xneg.txt",net0.n_1_2_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_5_ypos.txt",net0.n_1_2_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_5_yneg.txt",net0.n_1_2_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_5_zpos.txt",net0.n_1_2_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_5_zneg.txt",net0.n_1_2_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_5_xpos.txt",net0.n_1_2_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_5_xneg.txt",net0.n_1_2_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_5_ypos.txt",net0.n_1_2_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_5_yneg.txt",net0.n_1_2_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_5_zpos.txt",net0.n_1_2_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_5_zneg.txt",net0.n_1_2_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_5_xpos.txt",net0.n_1_2_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_5_xneg.txt",net0.n_1_2_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_5_ypos.txt",net0.n_1_2_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_5_yneg.txt",net0.n_1_2_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_5_zpos.txt",net0.n_1_2_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_5_zneg.txt",net0.n_1_2_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_6_local.txt",net0.n_1_2_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_6_xpos.txt",net0.n_1_2_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_6_xneg.txt",net0.n_1_2_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_6_ypos.txt",net0.n_1_2_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_6_yneg.txt",net0.n_1_2_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_6_zpos.txt",net0.n_1_2_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_6_zneg.txt",net0.n_1_2_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_6_xpos.txt",net0.n_1_2_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_6_xneg.txt",net0.n_1_2_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_6_ypos.txt",net0.n_1_2_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_6_yneg.txt",net0.n_1_2_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_6_zpos.txt",net0.n_1_2_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_6_zneg.txt",net0.n_1_2_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_6_xpos.txt",net0.n_1_2_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_6_xneg.txt",net0.n_1_2_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_6_ypos.txt",net0.n_1_2_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_6_yneg.txt",net0.n_1_2_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_6_zpos.txt",net0.n_1_2_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_6_zneg.txt",net0.n_1_2_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_7_local.txt",net0.n_1_2_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_7_xpos.txt",net0.n_1_2_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_7_xneg.txt",net0.n_1_2_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_7_ypos.txt",net0.n_1_2_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_7_yneg.txt",net0.n_1_2_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_7_zpos.txt",net0.n_1_2_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_2_7_zneg.txt",net0.n_1_2_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_7_xpos.txt",net0.n_1_2_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_7_xneg.txt",net0.n_1_2_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_7_ypos.txt",net0.n_1_2_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_7_yneg.txt",net0.n_1_2_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_7_zpos.txt",net0.n_1_2_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_2_7_zneg.txt",net0.n_1_2_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_7_xpos.txt",net0.n_1_2_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_7_xneg.txt",net0.n_1_2_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_7_ypos.txt",net0.n_1_2_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_7_yneg.txt",net0.n_1_2_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_7_zpos.txt",net0.n_1_2_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_2_7_zneg.txt",net0.n_1_2_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_0_local.txt",net0.n_1_3_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_0_xpos.txt",net0.n_1_3_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_0_xneg.txt",net0.n_1_3_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_0_ypos.txt",net0.n_1_3_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_0_yneg.txt",net0.n_1_3_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_0_zpos.txt",net0.n_1_3_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_0_zneg.txt",net0.n_1_3_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_0_xpos.txt",net0.n_1_3_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_0_xneg.txt",net0.n_1_3_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_0_ypos.txt",net0.n_1_3_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_0_yneg.txt",net0.n_1_3_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_0_zpos.txt",net0.n_1_3_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_0_zneg.txt",net0.n_1_3_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_0_xpos.txt",net0.n_1_3_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_0_xneg.txt",net0.n_1_3_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_0_ypos.txt",net0.n_1_3_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_0_yneg.txt",net0.n_1_3_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_0_zpos.txt",net0.n_1_3_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_0_zneg.txt",net0.n_1_3_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_1_local.txt",net0.n_1_3_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_1_xpos.txt",net0.n_1_3_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_1_xneg.txt",net0.n_1_3_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_1_ypos.txt",net0.n_1_3_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_1_yneg.txt",net0.n_1_3_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_1_zpos.txt",net0.n_1_3_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_1_zneg.txt",net0.n_1_3_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_1_xpos.txt",net0.n_1_3_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_1_xneg.txt",net0.n_1_3_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_1_ypos.txt",net0.n_1_3_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_1_yneg.txt",net0.n_1_3_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_1_zpos.txt",net0.n_1_3_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_1_zneg.txt",net0.n_1_3_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_1_xpos.txt",net0.n_1_3_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_1_xneg.txt",net0.n_1_3_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_1_ypos.txt",net0.n_1_3_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_1_yneg.txt",net0.n_1_3_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_1_zpos.txt",net0.n_1_3_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_1_zneg.txt",net0.n_1_3_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_2_local.txt",net0.n_1_3_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_2_xpos.txt",net0.n_1_3_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_2_xneg.txt",net0.n_1_3_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_2_ypos.txt",net0.n_1_3_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_2_yneg.txt",net0.n_1_3_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_2_zpos.txt",net0.n_1_3_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_2_zneg.txt",net0.n_1_3_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_2_xpos.txt",net0.n_1_3_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_2_xneg.txt",net0.n_1_3_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_2_ypos.txt",net0.n_1_3_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_2_yneg.txt",net0.n_1_3_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_2_zpos.txt",net0.n_1_3_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_2_zneg.txt",net0.n_1_3_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_2_xpos.txt",net0.n_1_3_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_2_xneg.txt",net0.n_1_3_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_2_ypos.txt",net0.n_1_3_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_2_yneg.txt",net0.n_1_3_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_2_zpos.txt",net0.n_1_3_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_2_zneg.txt",net0.n_1_3_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_3_local.txt",net0.n_1_3_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_3_xpos.txt",net0.n_1_3_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_3_xneg.txt",net0.n_1_3_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_3_ypos.txt",net0.n_1_3_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_3_yneg.txt",net0.n_1_3_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_3_zpos.txt",net0.n_1_3_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_3_zneg.txt",net0.n_1_3_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_3_xpos.txt",net0.n_1_3_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_3_xneg.txt",net0.n_1_3_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_3_ypos.txt",net0.n_1_3_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_3_yneg.txt",net0.n_1_3_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_3_zpos.txt",net0.n_1_3_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_3_zneg.txt",net0.n_1_3_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_3_xpos.txt",net0.n_1_3_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_3_xneg.txt",net0.n_1_3_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_3_ypos.txt",net0.n_1_3_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_3_yneg.txt",net0.n_1_3_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_3_zpos.txt",net0.n_1_3_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_3_zneg.txt",net0.n_1_3_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_4_local.txt",net0.n_1_3_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_4_xpos.txt",net0.n_1_3_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_4_xneg.txt",net0.n_1_3_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_4_ypos.txt",net0.n_1_3_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_4_yneg.txt",net0.n_1_3_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_4_zpos.txt",net0.n_1_3_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_4_zneg.txt",net0.n_1_3_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_4_xpos.txt",net0.n_1_3_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_4_xneg.txt",net0.n_1_3_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_4_ypos.txt",net0.n_1_3_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_4_yneg.txt",net0.n_1_3_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_4_zpos.txt",net0.n_1_3_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_4_zneg.txt",net0.n_1_3_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_4_xpos.txt",net0.n_1_3_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_4_xneg.txt",net0.n_1_3_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_4_ypos.txt",net0.n_1_3_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_4_yneg.txt",net0.n_1_3_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_4_zpos.txt",net0.n_1_3_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_4_zneg.txt",net0.n_1_3_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_5_local.txt",net0.n_1_3_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_5_xpos.txt",net0.n_1_3_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_5_xneg.txt",net0.n_1_3_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_5_ypos.txt",net0.n_1_3_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_5_yneg.txt",net0.n_1_3_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_5_zpos.txt",net0.n_1_3_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_5_zneg.txt",net0.n_1_3_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_5_xpos.txt",net0.n_1_3_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_5_xneg.txt",net0.n_1_3_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_5_ypos.txt",net0.n_1_3_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_5_yneg.txt",net0.n_1_3_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_5_zpos.txt",net0.n_1_3_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_5_zneg.txt",net0.n_1_3_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_5_xpos.txt",net0.n_1_3_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_5_xneg.txt",net0.n_1_3_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_5_ypos.txt",net0.n_1_3_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_5_yneg.txt",net0.n_1_3_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_5_zpos.txt",net0.n_1_3_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_5_zneg.txt",net0.n_1_3_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_6_local.txt",net0.n_1_3_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_6_xpos.txt",net0.n_1_3_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_6_xneg.txt",net0.n_1_3_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_6_ypos.txt",net0.n_1_3_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_6_yneg.txt",net0.n_1_3_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_6_zpos.txt",net0.n_1_3_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_6_zneg.txt",net0.n_1_3_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_6_xpos.txt",net0.n_1_3_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_6_xneg.txt",net0.n_1_3_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_6_ypos.txt",net0.n_1_3_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_6_yneg.txt",net0.n_1_3_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_6_zpos.txt",net0.n_1_3_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_6_zneg.txt",net0.n_1_3_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_6_xpos.txt",net0.n_1_3_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_6_xneg.txt",net0.n_1_3_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_6_ypos.txt",net0.n_1_3_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_6_yneg.txt",net0.n_1_3_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_6_zpos.txt",net0.n_1_3_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_6_zneg.txt",net0.n_1_3_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_7_local.txt",net0.n_1_3_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_7_xpos.txt",net0.n_1_3_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_7_xneg.txt",net0.n_1_3_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_7_ypos.txt",net0.n_1_3_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_7_yneg.txt",net0.n_1_3_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_7_zpos.txt",net0.n_1_3_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_3_7_zneg.txt",net0.n_1_3_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_7_xpos.txt",net0.n_1_3_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_7_xneg.txt",net0.n_1_3_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_7_ypos.txt",net0.n_1_3_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_7_yneg.txt",net0.n_1_3_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_7_zpos.txt",net0.n_1_3_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_3_7_zneg.txt",net0.n_1_3_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_7_xpos.txt",net0.n_1_3_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_7_xneg.txt",net0.n_1_3_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_7_ypos.txt",net0.n_1_3_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_7_yneg.txt",net0.n_1_3_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_7_zpos.txt",net0.n_1_3_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_3_7_zneg.txt",net0.n_1_3_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_0_local.txt",net0.n_1_4_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_0_xpos.txt",net0.n_1_4_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_0_xneg.txt",net0.n_1_4_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_0_ypos.txt",net0.n_1_4_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_0_yneg.txt",net0.n_1_4_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_0_zpos.txt",net0.n_1_4_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_0_zneg.txt",net0.n_1_4_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_0_xpos.txt",net0.n_1_4_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_0_xneg.txt",net0.n_1_4_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_0_ypos.txt",net0.n_1_4_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_0_yneg.txt",net0.n_1_4_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_0_zpos.txt",net0.n_1_4_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_0_zneg.txt",net0.n_1_4_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_0_xpos.txt",net0.n_1_4_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_0_xneg.txt",net0.n_1_4_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_0_ypos.txt",net0.n_1_4_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_0_yneg.txt",net0.n_1_4_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_0_zpos.txt",net0.n_1_4_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_0_zneg.txt",net0.n_1_4_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_1_local.txt",net0.n_1_4_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_1_xpos.txt",net0.n_1_4_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_1_xneg.txt",net0.n_1_4_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_1_ypos.txt",net0.n_1_4_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_1_yneg.txt",net0.n_1_4_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_1_zpos.txt",net0.n_1_4_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_1_zneg.txt",net0.n_1_4_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_1_xpos.txt",net0.n_1_4_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_1_xneg.txt",net0.n_1_4_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_1_ypos.txt",net0.n_1_4_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_1_yneg.txt",net0.n_1_4_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_1_zpos.txt",net0.n_1_4_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_1_zneg.txt",net0.n_1_4_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_1_xpos.txt",net0.n_1_4_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_1_xneg.txt",net0.n_1_4_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_1_ypos.txt",net0.n_1_4_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_1_yneg.txt",net0.n_1_4_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_1_zpos.txt",net0.n_1_4_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_1_zneg.txt",net0.n_1_4_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_2_local.txt",net0.n_1_4_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_2_xpos.txt",net0.n_1_4_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_2_xneg.txt",net0.n_1_4_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_2_ypos.txt",net0.n_1_4_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_2_yneg.txt",net0.n_1_4_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_2_zpos.txt",net0.n_1_4_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_2_zneg.txt",net0.n_1_4_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_2_xpos.txt",net0.n_1_4_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_2_xneg.txt",net0.n_1_4_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_2_ypos.txt",net0.n_1_4_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_2_yneg.txt",net0.n_1_4_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_2_zpos.txt",net0.n_1_4_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_2_zneg.txt",net0.n_1_4_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_2_xpos.txt",net0.n_1_4_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_2_xneg.txt",net0.n_1_4_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_2_ypos.txt",net0.n_1_4_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_2_yneg.txt",net0.n_1_4_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_2_zpos.txt",net0.n_1_4_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_2_zneg.txt",net0.n_1_4_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_3_local.txt",net0.n_1_4_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_3_xpos.txt",net0.n_1_4_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_3_xneg.txt",net0.n_1_4_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_3_ypos.txt",net0.n_1_4_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_3_yneg.txt",net0.n_1_4_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_3_zpos.txt",net0.n_1_4_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_3_zneg.txt",net0.n_1_4_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_3_xpos.txt",net0.n_1_4_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_3_xneg.txt",net0.n_1_4_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_3_ypos.txt",net0.n_1_4_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_3_yneg.txt",net0.n_1_4_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_3_zpos.txt",net0.n_1_4_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_3_zneg.txt",net0.n_1_4_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_3_xpos.txt",net0.n_1_4_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_3_xneg.txt",net0.n_1_4_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_3_ypos.txt",net0.n_1_4_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_3_yneg.txt",net0.n_1_4_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_3_zpos.txt",net0.n_1_4_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_3_zneg.txt",net0.n_1_4_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_4_local.txt",net0.n_1_4_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_4_xpos.txt",net0.n_1_4_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_4_xneg.txt",net0.n_1_4_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_4_ypos.txt",net0.n_1_4_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_4_yneg.txt",net0.n_1_4_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_4_zpos.txt",net0.n_1_4_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_4_zneg.txt",net0.n_1_4_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_4_xpos.txt",net0.n_1_4_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_4_xneg.txt",net0.n_1_4_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_4_ypos.txt",net0.n_1_4_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_4_yneg.txt",net0.n_1_4_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_4_zpos.txt",net0.n_1_4_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_4_zneg.txt",net0.n_1_4_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_4_xpos.txt",net0.n_1_4_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_4_xneg.txt",net0.n_1_4_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_4_ypos.txt",net0.n_1_4_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_4_yneg.txt",net0.n_1_4_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_4_zpos.txt",net0.n_1_4_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_4_zneg.txt",net0.n_1_4_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_5_local.txt",net0.n_1_4_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_5_xpos.txt",net0.n_1_4_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_5_xneg.txt",net0.n_1_4_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_5_ypos.txt",net0.n_1_4_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_5_yneg.txt",net0.n_1_4_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_5_zpos.txt",net0.n_1_4_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_5_zneg.txt",net0.n_1_4_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_5_xpos.txt",net0.n_1_4_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_5_xneg.txt",net0.n_1_4_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_5_ypos.txt",net0.n_1_4_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_5_yneg.txt",net0.n_1_4_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_5_zpos.txt",net0.n_1_4_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_5_zneg.txt",net0.n_1_4_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_5_xpos.txt",net0.n_1_4_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_5_xneg.txt",net0.n_1_4_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_5_ypos.txt",net0.n_1_4_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_5_yneg.txt",net0.n_1_4_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_5_zpos.txt",net0.n_1_4_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_5_zneg.txt",net0.n_1_4_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_6_local.txt",net0.n_1_4_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_6_xpos.txt",net0.n_1_4_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_6_xneg.txt",net0.n_1_4_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_6_ypos.txt",net0.n_1_4_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_6_yneg.txt",net0.n_1_4_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_6_zpos.txt",net0.n_1_4_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_6_zneg.txt",net0.n_1_4_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_6_xpos.txt",net0.n_1_4_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_6_xneg.txt",net0.n_1_4_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_6_ypos.txt",net0.n_1_4_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_6_yneg.txt",net0.n_1_4_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_6_zpos.txt",net0.n_1_4_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_6_zneg.txt",net0.n_1_4_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_6_xpos.txt",net0.n_1_4_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_6_xneg.txt",net0.n_1_4_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_6_ypos.txt",net0.n_1_4_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_6_yneg.txt",net0.n_1_4_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_6_zpos.txt",net0.n_1_4_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_6_zneg.txt",net0.n_1_4_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_7_local.txt",net0.n_1_4_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_7_xpos.txt",net0.n_1_4_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_7_xneg.txt",net0.n_1_4_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_7_ypos.txt",net0.n_1_4_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_7_yneg.txt",net0.n_1_4_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_7_zpos.txt",net0.n_1_4_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_4_7_zneg.txt",net0.n_1_4_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_7_xpos.txt",net0.n_1_4_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_7_xneg.txt",net0.n_1_4_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_7_ypos.txt",net0.n_1_4_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_7_yneg.txt",net0.n_1_4_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_7_zpos.txt",net0.n_1_4_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_4_7_zneg.txt",net0.n_1_4_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_7_xpos.txt",net0.n_1_4_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_7_xneg.txt",net0.n_1_4_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_7_ypos.txt",net0.n_1_4_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_7_yneg.txt",net0.n_1_4_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_7_zpos.txt",net0.n_1_4_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_4_7_zneg.txt",net0.n_1_4_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_0_local.txt",net0.n_1_5_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_0_xpos.txt",net0.n_1_5_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_0_xneg.txt",net0.n_1_5_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_0_ypos.txt",net0.n_1_5_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_0_yneg.txt",net0.n_1_5_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_0_zpos.txt",net0.n_1_5_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_0_zneg.txt",net0.n_1_5_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_0_xpos.txt",net0.n_1_5_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_0_xneg.txt",net0.n_1_5_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_0_ypos.txt",net0.n_1_5_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_0_yneg.txt",net0.n_1_5_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_0_zpos.txt",net0.n_1_5_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_0_zneg.txt",net0.n_1_5_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_0_xpos.txt",net0.n_1_5_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_0_xneg.txt",net0.n_1_5_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_0_ypos.txt",net0.n_1_5_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_0_yneg.txt",net0.n_1_5_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_0_zpos.txt",net0.n_1_5_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_0_zneg.txt",net0.n_1_5_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_1_local.txt",net0.n_1_5_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_1_xpos.txt",net0.n_1_5_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_1_xneg.txt",net0.n_1_5_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_1_ypos.txt",net0.n_1_5_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_1_yneg.txt",net0.n_1_5_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_1_zpos.txt",net0.n_1_5_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_1_zneg.txt",net0.n_1_5_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_1_xpos.txt",net0.n_1_5_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_1_xneg.txt",net0.n_1_5_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_1_ypos.txt",net0.n_1_5_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_1_yneg.txt",net0.n_1_5_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_1_zpos.txt",net0.n_1_5_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_1_zneg.txt",net0.n_1_5_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_1_xpos.txt",net0.n_1_5_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_1_xneg.txt",net0.n_1_5_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_1_ypos.txt",net0.n_1_5_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_1_yneg.txt",net0.n_1_5_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_1_zpos.txt",net0.n_1_5_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_1_zneg.txt",net0.n_1_5_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_2_local.txt",net0.n_1_5_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_2_xpos.txt",net0.n_1_5_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_2_xneg.txt",net0.n_1_5_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_2_ypos.txt",net0.n_1_5_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_2_yneg.txt",net0.n_1_5_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_2_zpos.txt",net0.n_1_5_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_2_zneg.txt",net0.n_1_5_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_2_xpos.txt",net0.n_1_5_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_2_xneg.txt",net0.n_1_5_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_2_ypos.txt",net0.n_1_5_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_2_yneg.txt",net0.n_1_5_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_2_zpos.txt",net0.n_1_5_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_2_zneg.txt",net0.n_1_5_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_2_xpos.txt",net0.n_1_5_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_2_xneg.txt",net0.n_1_5_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_2_ypos.txt",net0.n_1_5_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_2_yneg.txt",net0.n_1_5_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_2_zpos.txt",net0.n_1_5_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_2_zneg.txt",net0.n_1_5_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_3_local.txt",net0.n_1_5_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_3_xpos.txt",net0.n_1_5_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_3_xneg.txt",net0.n_1_5_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_3_ypos.txt",net0.n_1_5_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_3_yneg.txt",net0.n_1_5_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_3_zpos.txt",net0.n_1_5_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_3_zneg.txt",net0.n_1_5_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_3_xpos.txt",net0.n_1_5_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_3_xneg.txt",net0.n_1_5_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_3_ypos.txt",net0.n_1_5_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_3_yneg.txt",net0.n_1_5_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_3_zpos.txt",net0.n_1_5_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_3_zneg.txt",net0.n_1_5_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_3_xpos.txt",net0.n_1_5_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_3_xneg.txt",net0.n_1_5_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_3_ypos.txt",net0.n_1_5_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_3_yneg.txt",net0.n_1_5_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_3_zpos.txt",net0.n_1_5_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_3_zneg.txt",net0.n_1_5_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_4_local.txt",net0.n_1_5_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_4_xpos.txt",net0.n_1_5_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_4_xneg.txt",net0.n_1_5_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_4_ypos.txt",net0.n_1_5_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_4_yneg.txt",net0.n_1_5_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_4_zpos.txt",net0.n_1_5_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_4_zneg.txt",net0.n_1_5_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_4_xpos.txt",net0.n_1_5_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_4_xneg.txt",net0.n_1_5_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_4_ypos.txt",net0.n_1_5_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_4_yneg.txt",net0.n_1_5_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_4_zpos.txt",net0.n_1_5_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_4_zneg.txt",net0.n_1_5_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_4_xpos.txt",net0.n_1_5_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_4_xneg.txt",net0.n_1_5_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_4_ypos.txt",net0.n_1_5_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_4_yneg.txt",net0.n_1_5_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_4_zpos.txt",net0.n_1_5_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_4_zneg.txt",net0.n_1_5_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_5_local.txt",net0.n_1_5_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_5_xpos.txt",net0.n_1_5_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_5_xneg.txt",net0.n_1_5_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_5_ypos.txt",net0.n_1_5_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_5_yneg.txt",net0.n_1_5_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_5_zpos.txt",net0.n_1_5_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_5_zneg.txt",net0.n_1_5_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_5_xpos.txt",net0.n_1_5_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_5_xneg.txt",net0.n_1_5_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_5_ypos.txt",net0.n_1_5_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_5_yneg.txt",net0.n_1_5_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_5_zpos.txt",net0.n_1_5_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_5_zneg.txt",net0.n_1_5_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_5_xpos.txt",net0.n_1_5_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_5_xneg.txt",net0.n_1_5_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_5_ypos.txt",net0.n_1_5_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_5_yneg.txt",net0.n_1_5_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_5_zpos.txt",net0.n_1_5_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_5_zneg.txt",net0.n_1_5_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_6_local.txt",net0.n_1_5_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_6_xpos.txt",net0.n_1_5_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_6_xneg.txt",net0.n_1_5_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_6_ypos.txt",net0.n_1_5_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_6_yneg.txt",net0.n_1_5_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_6_zpos.txt",net0.n_1_5_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_6_zneg.txt",net0.n_1_5_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_6_xpos.txt",net0.n_1_5_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_6_xneg.txt",net0.n_1_5_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_6_ypos.txt",net0.n_1_5_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_6_yneg.txt",net0.n_1_5_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_6_zpos.txt",net0.n_1_5_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_6_zneg.txt",net0.n_1_5_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_6_xpos.txt",net0.n_1_5_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_6_xneg.txt",net0.n_1_5_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_6_ypos.txt",net0.n_1_5_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_6_yneg.txt",net0.n_1_5_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_6_zpos.txt",net0.n_1_5_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_6_zneg.txt",net0.n_1_5_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_7_local.txt",net0.n_1_5_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_7_xpos.txt",net0.n_1_5_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_7_xneg.txt",net0.n_1_5_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_7_ypos.txt",net0.n_1_5_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_7_yneg.txt",net0.n_1_5_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_7_zpos.txt",net0.n_1_5_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_5_7_zneg.txt",net0.n_1_5_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_7_xpos.txt",net0.n_1_5_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_7_xneg.txt",net0.n_1_5_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_7_ypos.txt",net0.n_1_5_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_7_yneg.txt",net0.n_1_5_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_7_zpos.txt",net0.n_1_5_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_5_7_zneg.txt",net0.n_1_5_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_7_xpos.txt",net0.n_1_5_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_7_xneg.txt",net0.n_1_5_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_7_ypos.txt",net0.n_1_5_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_7_yneg.txt",net0.n_1_5_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_7_zpos.txt",net0.n_1_5_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_5_7_zneg.txt",net0.n_1_5_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_0_local.txt",net0.n_1_6_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_0_xpos.txt",net0.n_1_6_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_0_xneg.txt",net0.n_1_6_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_0_ypos.txt",net0.n_1_6_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_0_yneg.txt",net0.n_1_6_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_0_zpos.txt",net0.n_1_6_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_0_zneg.txt",net0.n_1_6_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_0_xpos.txt",net0.n_1_6_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_0_xneg.txt",net0.n_1_6_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_0_ypos.txt",net0.n_1_6_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_0_yneg.txt",net0.n_1_6_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_0_zpos.txt",net0.n_1_6_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_0_zneg.txt",net0.n_1_6_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_0_xpos.txt",net0.n_1_6_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_0_xneg.txt",net0.n_1_6_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_0_ypos.txt",net0.n_1_6_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_0_yneg.txt",net0.n_1_6_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_0_zpos.txt",net0.n_1_6_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_0_zneg.txt",net0.n_1_6_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_1_local.txt",net0.n_1_6_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_1_xpos.txt",net0.n_1_6_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_1_xneg.txt",net0.n_1_6_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_1_ypos.txt",net0.n_1_6_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_1_yneg.txt",net0.n_1_6_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_1_zpos.txt",net0.n_1_6_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_1_zneg.txt",net0.n_1_6_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_1_xpos.txt",net0.n_1_6_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_1_xneg.txt",net0.n_1_6_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_1_ypos.txt",net0.n_1_6_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_1_yneg.txt",net0.n_1_6_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_1_zpos.txt",net0.n_1_6_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_1_zneg.txt",net0.n_1_6_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_1_xpos.txt",net0.n_1_6_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_1_xneg.txt",net0.n_1_6_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_1_ypos.txt",net0.n_1_6_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_1_yneg.txt",net0.n_1_6_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_1_zpos.txt",net0.n_1_6_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_1_zneg.txt",net0.n_1_6_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_2_local.txt",net0.n_1_6_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_2_xpos.txt",net0.n_1_6_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_2_xneg.txt",net0.n_1_6_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_2_ypos.txt",net0.n_1_6_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_2_yneg.txt",net0.n_1_6_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_2_zpos.txt",net0.n_1_6_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_2_zneg.txt",net0.n_1_6_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_2_xpos.txt",net0.n_1_6_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_2_xneg.txt",net0.n_1_6_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_2_ypos.txt",net0.n_1_6_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_2_yneg.txt",net0.n_1_6_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_2_zpos.txt",net0.n_1_6_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_2_zneg.txt",net0.n_1_6_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_2_xpos.txt",net0.n_1_6_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_2_xneg.txt",net0.n_1_6_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_2_ypos.txt",net0.n_1_6_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_2_yneg.txt",net0.n_1_6_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_2_zpos.txt",net0.n_1_6_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_2_zneg.txt",net0.n_1_6_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_3_local.txt",net0.n_1_6_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_3_xpos.txt",net0.n_1_6_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_3_xneg.txt",net0.n_1_6_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_3_ypos.txt",net0.n_1_6_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_3_yneg.txt",net0.n_1_6_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_3_zpos.txt",net0.n_1_6_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_3_zneg.txt",net0.n_1_6_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_3_xpos.txt",net0.n_1_6_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_3_xneg.txt",net0.n_1_6_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_3_ypos.txt",net0.n_1_6_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_3_yneg.txt",net0.n_1_6_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_3_zpos.txt",net0.n_1_6_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_3_zneg.txt",net0.n_1_6_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_3_xpos.txt",net0.n_1_6_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_3_xneg.txt",net0.n_1_6_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_3_ypos.txt",net0.n_1_6_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_3_yneg.txt",net0.n_1_6_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_3_zpos.txt",net0.n_1_6_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_3_zneg.txt",net0.n_1_6_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_4_local.txt",net0.n_1_6_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_4_xpos.txt",net0.n_1_6_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_4_xneg.txt",net0.n_1_6_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_4_ypos.txt",net0.n_1_6_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_4_yneg.txt",net0.n_1_6_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_4_zpos.txt",net0.n_1_6_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_4_zneg.txt",net0.n_1_6_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_4_xpos.txt",net0.n_1_6_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_4_xneg.txt",net0.n_1_6_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_4_ypos.txt",net0.n_1_6_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_4_yneg.txt",net0.n_1_6_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_4_zpos.txt",net0.n_1_6_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_4_zneg.txt",net0.n_1_6_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_4_xpos.txt",net0.n_1_6_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_4_xneg.txt",net0.n_1_6_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_4_ypos.txt",net0.n_1_6_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_4_yneg.txt",net0.n_1_6_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_4_zpos.txt",net0.n_1_6_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_4_zneg.txt",net0.n_1_6_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_5_local.txt",net0.n_1_6_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_5_xpos.txt",net0.n_1_6_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_5_xneg.txt",net0.n_1_6_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_5_ypos.txt",net0.n_1_6_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_5_yneg.txt",net0.n_1_6_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_5_zpos.txt",net0.n_1_6_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_5_zneg.txt",net0.n_1_6_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_5_xpos.txt",net0.n_1_6_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_5_xneg.txt",net0.n_1_6_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_5_ypos.txt",net0.n_1_6_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_5_yneg.txt",net0.n_1_6_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_5_zpos.txt",net0.n_1_6_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_5_zneg.txt",net0.n_1_6_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_5_xpos.txt",net0.n_1_6_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_5_xneg.txt",net0.n_1_6_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_5_ypos.txt",net0.n_1_6_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_5_yneg.txt",net0.n_1_6_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_5_zpos.txt",net0.n_1_6_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_5_zneg.txt",net0.n_1_6_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_6_local.txt",net0.n_1_6_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_6_xpos.txt",net0.n_1_6_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_6_xneg.txt",net0.n_1_6_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_6_ypos.txt",net0.n_1_6_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_6_yneg.txt",net0.n_1_6_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_6_zpos.txt",net0.n_1_6_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_6_zneg.txt",net0.n_1_6_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_6_xpos.txt",net0.n_1_6_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_6_xneg.txt",net0.n_1_6_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_6_ypos.txt",net0.n_1_6_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_6_yneg.txt",net0.n_1_6_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_6_zpos.txt",net0.n_1_6_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_6_zneg.txt",net0.n_1_6_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_6_xpos.txt",net0.n_1_6_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_6_xneg.txt",net0.n_1_6_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_6_ypos.txt",net0.n_1_6_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_6_yneg.txt",net0.n_1_6_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_6_zpos.txt",net0.n_1_6_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_6_zneg.txt",net0.n_1_6_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_7_local.txt",net0.n_1_6_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_7_xpos.txt",net0.n_1_6_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_7_xneg.txt",net0.n_1_6_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_7_ypos.txt",net0.n_1_6_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_7_yneg.txt",net0.n_1_6_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_7_zpos.txt",net0.n_1_6_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_6_7_zneg.txt",net0.n_1_6_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_7_xpos.txt",net0.n_1_6_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_7_xneg.txt",net0.n_1_6_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_7_ypos.txt",net0.n_1_6_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_7_yneg.txt",net0.n_1_6_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_7_zpos.txt",net0.n_1_6_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_6_7_zneg.txt",net0.n_1_6_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_7_xpos.txt",net0.n_1_6_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_7_xneg.txt",net0.n_1_6_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_7_ypos.txt",net0.n_1_6_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_7_yneg.txt",net0.n_1_6_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_7_zpos.txt",net0.n_1_6_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_6_7_zneg.txt",net0.n_1_6_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_0_local.txt",net0.n_1_7_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_0_xpos.txt",net0.n_1_7_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_0_xneg.txt",net0.n_1_7_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_0_ypos.txt",net0.n_1_7_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_0_yneg.txt",net0.n_1_7_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_0_zpos.txt",net0.n_1_7_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_0_zneg.txt",net0.n_1_7_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_0_xpos.txt",net0.n_1_7_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_0_xneg.txt",net0.n_1_7_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_0_ypos.txt",net0.n_1_7_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_0_yneg.txt",net0.n_1_7_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_0_zpos.txt",net0.n_1_7_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_0_zneg.txt",net0.n_1_7_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_0_xpos.txt",net0.n_1_7_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_0_xneg.txt",net0.n_1_7_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_0_ypos.txt",net0.n_1_7_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_0_yneg.txt",net0.n_1_7_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_0_zpos.txt",net0.n_1_7_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_0_zneg.txt",net0.n_1_7_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_1_local.txt",net0.n_1_7_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_1_xpos.txt",net0.n_1_7_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_1_xneg.txt",net0.n_1_7_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_1_ypos.txt",net0.n_1_7_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_1_yneg.txt",net0.n_1_7_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_1_zpos.txt",net0.n_1_7_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_1_zneg.txt",net0.n_1_7_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_1_xpos.txt",net0.n_1_7_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_1_xneg.txt",net0.n_1_7_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_1_ypos.txt",net0.n_1_7_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_1_yneg.txt",net0.n_1_7_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_1_zpos.txt",net0.n_1_7_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_1_zneg.txt",net0.n_1_7_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_1_xpos.txt",net0.n_1_7_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_1_xneg.txt",net0.n_1_7_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_1_ypos.txt",net0.n_1_7_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_1_yneg.txt",net0.n_1_7_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_1_zpos.txt",net0.n_1_7_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_1_zneg.txt",net0.n_1_7_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_2_local.txt",net0.n_1_7_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_2_xpos.txt",net0.n_1_7_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_2_xneg.txt",net0.n_1_7_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_2_ypos.txt",net0.n_1_7_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_2_yneg.txt",net0.n_1_7_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_2_zpos.txt",net0.n_1_7_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_2_zneg.txt",net0.n_1_7_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_2_xpos.txt",net0.n_1_7_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_2_xneg.txt",net0.n_1_7_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_2_ypos.txt",net0.n_1_7_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_2_yneg.txt",net0.n_1_7_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_2_zpos.txt",net0.n_1_7_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_2_zneg.txt",net0.n_1_7_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_2_xpos.txt",net0.n_1_7_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_2_xneg.txt",net0.n_1_7_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_2_ypos.txt",net0.n_1_7_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_2_yneg.txt",net0.n_1_7_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_2_zpos.txt",net0.n_1_7_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_2_zneg.txt",net0.n_1_7_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_3_local.txt",net0.n_1_7_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_3_xpos.txt",net0.n_1_7_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_3_xneg.txt",net0.n_1_7_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_3_ypos.txt",net0.n_1_7_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_3_yneg.txt",net0.n_1_7_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_3_zpos.txt",net0.n_1_7_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_3_zneg.txt",net0.n_1_7_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_3_xpos.txt",net0.n_1_7_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_3_xneg.txt",net0.n_1_7_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_3_ypos.txt",net0.n_1_7_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_3_yneg.txt",net0.n_1_7_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_3_zpos.txt",net0.n_1_7_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_3_zneg.txt",net0.n_1_7_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_3_xpos.txt",net0.n_1_7_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_3_xneg.txt",net0.n_1_7_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_3_ypos.txt",net0.n_1_7_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_3_yneg.txt",net0.n_1_7_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_3_zpos.txt",net0.n_1_7_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_3_zneg.txt",net0.n_1_7_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_4_local.txt",net0.n_1_7_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_4_xpos.txt",net0.n_1_7_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_4_xneg.txt",net0.n_1_7_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_4_ypos.txt",net0.n_1_7_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_4_yneg.txt",net0.n_1_7_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_4_zpos.txt",net0.n_1_7_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_4_zneg.txt",net0.n_1_7_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_4_xpos.txt",net0.n_1_7_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_4_xneg.txt",net0.n_1_7_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_4_ypos.txt",net0.n_1_7_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_4_yneg.txt",net0.n_1_7_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_4_zpos.txt",net0.n_1_7_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_4_zneg.txt",net0.n_1_7_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_4_xpos.txt",net0.n_1_7_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_4_xneg.txt",net0.n_1_7_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_4_ypos.txt",net0.n_1_7_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_4_yneg.txt",net0.n_1_7_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_4_zpos.txt",net0.n_1_7_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_4_zneg.txt",net0.n_1_7_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_5_local.txt",net0.n_1_7_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_5_xpos.txt",net0.n_1_7_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_5_xneg.txt",net0.n_1_7_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_5_ypos.txt",net0.n_1_7_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_5_yneg.txt",net0.n_1_7_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_5_zpos.txt",net0.n_1_7_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_5_zneg.txt",net0.n_1_7_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_5_xpos.txt",net0.n_1_7_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_5_xneg.txt",net0.n_1_7_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_5_ypos.txt",net0.n_1_7_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_5_yneg.txt",net0.n_1_7_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_5_zpos.txt",net0.n_1_7_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_5_zneg.txt",net0.n_1_7_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_5_xpos.txt",net0.n_1_7_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_5_xneg.txt",net0.n_1_7_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_5_ypos.txt",net0.n_1_7_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_5_yneg.txt",net0.n_1_7_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_5_zpos.txt",net0.n_1_7_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_5_zneg.txt",net0.n_1_7_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_6_local.txt",net0.n_1_7_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_6_xpos.txt",net0.n_1_7_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_6_xneg.txt",net0.n_1_7_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_6_ypos.txt",net0.n_1_7_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_6_yneg.txt",net0.n_1_7_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_6_zpos.txt",net0.n_1_7_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_6_zneg.txt",net0.n_1_7_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_6_xpos.txt",net0.n_1_7_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_6_xneg.txt",net0.n_1_7_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_6_ypos.txt",net0.n_1_7_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_6_yneg.txt",net0.n_1_7_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_6_zpos.txt",net0.n_1_7_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_6_zneg.txt",net0.n_1_7_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_6_xpos.txt",net0.n_1_7_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_6_xneg.txt",net0.n_1_7_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_6_ypos.txt",net0.n_1_7_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_6_yneg.txt",net0.n_1_7_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_6_zpos.txt",net0.n_1_7_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_6_zneg.txt",net0.n_1_7_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_7_local.txt",net0.n_1_7_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_7_xpos.txt",net0.n_1_7_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_7_xneg.txt",net0.n_1_7_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_7_ypos.txt",net0.n_1_7_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_7_yneg.txt",net0.n_1_7_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_7_zpos.txt",net0.n_1_7_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_1_7_7_zneg.txt",net0.n_1_7_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_7_xpos.txt",net0.n_1_7_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_7_xneg.txt",net0.n_1_7_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_7_ypos.txt",net0.n_1_7_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_7_yneg.txt",net0.n_1_7_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_7_zpos.txt",net0.n_1_7_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_1_7_7_zneg.txt",net0.n_1_7_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_7_xpos.txt",net0.n_1_7_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_7_xneg.txt",net0.n_1_7_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_7_ypos.txt",net0.n_1_7_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_7_yneg.txt",net0.n_1_7_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_7_zpos.txt",net0.n_1_7_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_1_7_7_zneg.txt",net0.n_1_7_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_0_local.txt",net0.n_2_0_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_0_xpos.txt",net0.n_2_0_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_0_xneg.txt",net0.n_2_0_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_0_ypos.txt",net0.n_2_0_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_0_yneg.txt",net0.n_2_0_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_0_zpos.txt",net0.n_2_0_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_0_zneg.txt",net0.n_2_0_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_0_xpos.txt",net0.n_2_0_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_0_xneg.txt",net0.n_2_0_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_0_ypos.txt",net0.n_2_0_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_0_yneg.txt",net0.n_2_0_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_0_zpos.txt",net0.n_2_0_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_0_zneg.txt",net0.n_2_0_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_0_xpos.txt",net0.n_2_0_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_0_xneg.txt",net0.n_2_0_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_0_ypos.txt",net0.n_2_0_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_0_yneg.txt",net0.n_2_0_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_0_zpos.txt",net0.n_2_0_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_0_zneg.txt",net0.n_2_0_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_1_local.txt",net0.n_2_0_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_1_xpos.txt",net0.n_2_0_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_1_xneg.txt",net0.n_2_0_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_1_ypos.txt",net0.n_2_0_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_1_yneg.txt",net0.n_2_0_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_1_zpos.txt",net0.n_2_0_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_1_zneg.txt",net0.n_2_0_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_1_xpos.txt",net0.n_2_0_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_1_xneg.txt",net0.n_2_0_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_1_ypos.txt",net0.n_2_0_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_1_yneg.txt",net0.n_2_0_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_1_zpos.txt",net0.n_2_0_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_1_zneg.txt",net0.n_2_0_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_1_xpos.txt",net0.n_2_0_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_1_xneg.txt",net0.n_2_0_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_1_ypos.txt",net0.n_2_0_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_1_yneg.txt",net0.n_2_0_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_1_zpos.txt",net0.n_2_0_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_1_zneg.txt",net0.n_2_0_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_2_local.txt",net0.n_2_0_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_2_xpos.txt",net0.n_2_0_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_2_xneg.txt",net0.n_2_0_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_2_ypos.txt",net0.n_2_0_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_2_yneg.txt",net0.n_2_0_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_2_zpos.txt",net0.n_2_0_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_2_zneg.txt",net0.n_2_0_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_2_xpos.txt",net0.n_2_0_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_2_xneg.txt",net0.n_2_0_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_2_ypos.txt",net0.n_2_0_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_2_yneg.txt",net0.n_2_0_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_2_zpos.txt",net0.n_2_0_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_2_zneg.txt",net0.n_2_0_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_2_xpos.txt",net0.n_2_0_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_2_xneg.txt",net0.n_2_0_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_2_ypos.txt",net0.n_2_0_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_2_yneg.txt",net0.n_2_0_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_2_zpos.txt",net0.n_2_0_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_2_zneg.txt",net0.n_2_0_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_3_local.txt",net0.n_2_0_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_3_xpos.txt",net0.n_2_0_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_3_xneg.txt",net0.n_2_0_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_3_ypos.txt",net0.n_2_0_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_3_yneg.txt",net0.n_2_0_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_3_zpos.txt",net0.n_2_0_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_3_zneg.txt",net0.n_2_0_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_3_xpos.txt",net0.n_2_0_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_3_xneg.txt",net0.n_2_0_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_3_ypos.txt",net0.n_2_0_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_3_yneg.txt",net0.n_2_0_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_3_zpos.txt",net0.n_2_0_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_3_zneg.txt",net0.n_2_0_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_3_xpos.txt",net0.n_2_0_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_3_xneg.txt",net0.n_2_0_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_3_ypos.txt",net0.n_2_0_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_3_yneg.txt",net0.n_2_0_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_3_zpos.txt",net0.n_2_0_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_3_zneg.txt",net0.n_2_0_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_4_local.txt",net0.n_2_0_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_4_xpos.txt",net0.n_2_0_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_4_xneg.txt",net0.n_2_0_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_4_ypos.txt",net0.n_2_0_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_4_yneg.txt",net0.n_2_0_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_4_zpos.txt",net0.n_2_0_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_4_zneg.txt",net0.n_2_0_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_4_xpos.txt",net0.n_2_0_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_4_xneg.txt",net0.n_2_0_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_4_ypos.txt",net0.n_2_0_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_4_yneg.txt",net0.n_2_0_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_4_zpos.txt",net0.n_2_0_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_4_zneg.txt",net0.n_2_0_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_4_xpos.txt",net0.n_2_0_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_4_xneg.txt",net0.n_2_0_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_4_ypos.txt",net0.n_2_0_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_4_yneg.txt",net0.n_2_0_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_4_zpos.txt",net0.n_2_0_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_4_zneg.txt",net0.n_2_0_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_5_local.txt",net0.n_2_0_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_5_xpos.txt",net0.n_2_0_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_5_xneg.txt",net0.n_2_0_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_5_ypos.txt",net0.n_2_0_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_5_yneg.txt",net0.n_2_0_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_5_zpos.txt",net0.n_2_0_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_5_zneg.txt",net0.n_2_0_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_5_xpos.txt",net0.n_2_0_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_5_xneg.txt",net0.n_2_0_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_5_ypos.txt",net0.n_2_0_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_5_yneg.txt",net0.n_2_0_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_5_zpos.txt",net0.n_2_0_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_5_zneg.txt",net0.n_2_0_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_5_xpos.txt",net0.n_2_0_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_5_xneg.txt",net0.n_2_0_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_5_ypos.txt",net0.n_2_0_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_5_yneg.txt",net0.n_2_0_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_5_zpos.txt",net0.n_2_0_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_5_zneg.txt",net0.n_2_0_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_6_local.txt",net0.n_2_0_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_6_xpos.txt",net0.n_2_0_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_6_xneg.txt",net0.n_2_0_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_6_ypos.txt",net0.n_2_0_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_6_yneg.txt",net0.n_2_0_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_6_zpos.txt",net0.n_2_0_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_6_zneg.txt",net0.n_2_0_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_6_xpos.txt",net0.n_2_0_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_6_xneg.txt",net0.n_2_0_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_6_ypos.txt",net0.n_2_0_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_6_yneg.txt",net0.n_2_0_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_6_zpos.txt",net0.n_2_0_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_6_zneg.txt",net0.n_2_0_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_6_xpos.txt",net0.n_2_0_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_6_xneg.txt",net0.n_2_0_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_6_ypos.txt",net0.n_2_0_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_6_yneg.txt",net0.n_2_0_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_6_zpos.txt",net0.n_2_0_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_6_zneg.txt",net0.n_2_0_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_7_local.txt",net0.n_2_0_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_7_xpos.txt",net0.n_2_0_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_7_xneg.txt",net0.n_2_0_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_7_ypos.txt",net0.n_2_0_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_7_yneg.txt",net0.n_2_0_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_7_zpos.txt",net0.n_2_0_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_0_7_zneg.txt",net0.n_2_0_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_7_xpos.txt",net0.n_2_0_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_7_xneg.txt",net0.n_2_0_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_7_ypos.txt",net0.n_2_0_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_7_yneg.txt",net0.n_2_0_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_7_zpos.txt",net0.n_2_0_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_0_7_zneg.txt",net0.n_2_0_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_7_xpos.txt",net0.n_2_0_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_7_xneg.txt",net0.n_2_0_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_7_ypos.txt",net0.n_2_0_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_7_yneg.txt",net0.n_2_0_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_7_zpos.txt",net0.n_2_0_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_0_7_zneg.txt",net0.n_2_0_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_0_local.txt",net0.n_2_1_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_0_xpos.txt",net0.n_2_1_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_0_xneg.txt",net0.n_2_1_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_0_ypos.txt",net0.n_2_1_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_0_yneg.txt",net0.n_2_1_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_0_zpos.txt",net0.n_2_1_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_0_zneg.txt",net0.n_2_1_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_0_xpos.txt",net0.n_2_1_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_0_xneg.txt",net0.n_2_1_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_0_ypos.txt",net0.n_2_1_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_0_yneg.txt",net0.n_2_1_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_0_zpos.txt",net0.n_2_1_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_0_zneg.txt",net0.n_2_1_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_0_xpos.txt",net0.n_2_1_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_0_xneg.txt",net0.n_2_1_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_0_ypos.txt",net0.n_2_1_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_0_yneg.txt",net0.n_2_1_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_0_zpos.txt",net0.n_2_1_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_0_zneg.txt",net0.n_2_1_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_1_local.txt",net0.n_2_1_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_1_xpos.txt",net0.n_2_1_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_1_xneg.txt",net0.n_2_1_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_1_ypos.txt",net0.n_2_1_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_1_yneg.txt",net0.n_2_1_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_1_zpos.txt",net0.n_2_1_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_1_zneg.txt",net0.n_2_1_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_1_xpos.txt",net0.n_2_1_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_1_xneg.txt",net0.n_2_1_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_1_ypos.txt",net0.n_2_1_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_1_yneg.txt",net0.n_2_1_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_1_zpos.txt",net0.n_2_1_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_1_zneg.txt",net0.n_2_1_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_1_xpos.txt",net0.n_2_1_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_1_xneg.txt",net0.n_2_1_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_1_ypos.txt",net0.n_2_1_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_1_yneg.txt",net0.n_2_1_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_1_zpos.txt",net0.n_2_1_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_1_zneg.txt",net0.n_2_1_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_2_local.txt",net0.n_2_1_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_2_xpos.txt",net0.n_2_1_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_2_xneg.txt",net0.n_2_1_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_2_ypos.txt",net0.n_2_1_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_2_yneg.txt",net0.n_2_1_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_2_zpos.txt",net0.n_2_1_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_2_zneg.txt",net0.n_2_1_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_2_xpos.txt",net0.n_2_1_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_2_xneg.txt",net0.n_2_1_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_2_ypos.txt",net0.n_2_1_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_2_yneg.txt",net0.n_2_1_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_2_zpos.txt",net0.n_2_1_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_2_zneg.txt",net0.n_2_1_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_2_xpos.txt",net0.n_2_1_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_2_xneg.txt",net0.n_2_1_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_2_ypos.txt",net0.n_2_1_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_2_yneg.txt",net0.n_2_1_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_2_zpos.txt",net0.n_2_1_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_2_zneg.txt",net0.n_2_1_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_3_local.txt",net0.n_2_1_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_3_xpos.txt",net0.n_2_1_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_3_xneg.txt",net0.n_2_1_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_3_ypos.txt",net0.n_2_1_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_3_yneg.txt",net0.n_2_1_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_3_zpos.txt",net0.n_2_1_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_3_zneg.txt",net0.n_2_1_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_3_xpos.txt",net0.n_2_1_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_3_xneg.txt",net0.n_2_1_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_3_ypos.txt",net0.n_2_1_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_3_yneg.txt",net0.n_2_1_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_3_zpos.txt",net0.n_2_1_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_3_zneg.txt",net0.n_2_1_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_3_xpos.txt",net0.n_2_1_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_3_xneg.txt",net0.n_2_1_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_3_ypos.txt",net0.n_2_1_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_3_yneg.txt",net0.n_2_1_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_3_zpos.txt",net0.n_2_1_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_3_zneg.txt",net0.n_2_1_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_4_local.txt",net0.n_2_1_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_4_xpos.txt",net0.n_2_1_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_4_xneg.txt",net0.n_2_1_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_4_ypos.txt",net0.n_2_1_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_4_yneg.txt",net0.n_2_1_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_4_zpos.txt",net0.n_2_1_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_4_zneg.txt",net0.n_2_1_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_4_xpos.txt",net0.n_2_1_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_4_xneg.txt",net0.n_2_1_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_4_ypos.txt",net0.n_2_1_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_4_yneg.txt",net0.n_2_1_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_4_zpos.txt",net0.n_2_1_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_4_zneg.txt",net0.n_2_1_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_4_xpos.txt",net0.n_2_1_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_4_xneg.txt",net0.n_2_1_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_4_ypos.txt",net0.n_2_1_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_4_yneg.txt",net0.n_2_1_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_4_zpos.txt",net0.n_2_1_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_4_zneg.txt",net0.n_2_1_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_5_local.txt",net0.n_2_1_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_5_xpos.txt",net0.n_2_1_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_5_xneg.txt",net0.n_2_1_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_5_ypos.txt",net0.n_2_1_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_5_yneg.txt",net0.n_2_1_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_5_zpos.txt",net0.n_2_1_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_5_zneg.txt",net0.n_2_1_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_5_xpos.txt",net0.n_2_1_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_5_xneg.txt",net0.n_2_1_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_5_ypos.txt",net0.n_2_1_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_5_yneg.txt",net0.n_2_1_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_5_zpos.txt",net0.n_2_1_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_5_zneg.txt",net0.n_2_1_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_5_xpos.txt",net0.n_2_1_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_5_xneg.txt",net0.n_2_1_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_5_ypos.txt",net0.n_2_1_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_5_yneg.txt",net0.n_2_1_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_5_zpos.txt",net0.n_2_1_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_5_zneg.txt",net0.n_2_1_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_6_local.txt",net0.n_2_1_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_6_xpos.txt",net0.n_2_1_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_6_xneg.txt",net0.n_2_1_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_6_ypos.txt",net0.n_2_1_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_6_yneg.txt",net0.n_2_1_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_6_zpos.txt",net0.n_2_1_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_6_zneg.txt",net0.n_2_1_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_6_xpos.txt",net0.n_2_1_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_6_xneg.txt",net0.n_2_1_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_6_ypos.txt",net0.n_2_1_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_6_yneg.txt",net0.n_2_1_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_6_zpos.txt",net0.n_2_1_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_6_zneg.txt",net0.n_2_1_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_6_xpos.txt",net0.n_2_1_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_6_xneg.txt",net0.n_2_1_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_6_ypos.txt",net0.n_2_1_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_6_yneg.txt",net0.n_2_1_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_6_zpos.txt",net0.n_2_1_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_6_zneg.txt",net0.n_2_1_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_7_local.txt",net0.n_2_1_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_7_xpos.txt",net0.n_2_1_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_7_xneg.txt",net0.n_2_1_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_7_ypos.txt",net0.n_2_1_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_7_yneg.txt",net0.n_2_1_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_7_zpos.txt",net0.n_2_1_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_1_7_zneg.txt",net0.n_2_1_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_7_xpos.txt",net0.n_2_1_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_7_xneg.txt",net0.n_2_1_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_7_ypos.txt",net0.n_2_1_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_7_yneg.txt",net0.n_2_1_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_7_zpos.txt",net0.n_2_1_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_1_7_zneg.txt",net0.n_2_1_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_7_xpos.txt",net0.n_2_1_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_7_xneg.txt",net0.n_2_1_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_7_ypos.txt",net0.n_2_1_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_7_yneg.txt",net0.n_2_1_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_7_zpos.txt",net0.n_2_1_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_1_7_zneg.txt",net0.n_2_1_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_0_local.txt",net0.n_2_2_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_0_xpos.txt",net0.n_2_2_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_0_xneg.txt",net0.n_2_2_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_0_ypos.txt",net0.n_2_2_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_0_yneg.txt",net0.n_2_2_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_0_zpos.txt",net0.n_2_2_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_0_zneg.txt",net0.n_2_2_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_0_xpos.txt",net0.n_2_2_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_0_xneg.txt",net0.n_2_2_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_0_ypos.txt",net0.n_2_2_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_0_yneg.txt",net0.n_2_2_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_0_zpos.txt",net0.n_2_2_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_0_zneg.txt",net0.n_2_2_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_0_xpos.txt",net0.n_2_2_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_0_xneg.txt",net0.n_2_2_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_0_ypos.txt",net0.n_2_2_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_0_yneg.txt",net0.n_2_2_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_0_zpos.txt",net0.n_2_2_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_0_zneg.txt",net0.n_2_2_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_1_local.txt",net0.n_2_2_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_1_xpos.txt",net0.n_2_2_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_1_xneg.txt",net0.n_2_2_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_1_ypos.txt",net0.n_2_2_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_1_yneg.txt",net0.n_2_2_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_1_zpos.txt",net0.n_2_2_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_1_zneg.txt",net0.n_2_2_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_1_xpos.txt",net0.n_2_2_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_1_xneg.txt",net0.n_2_2_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_1_ypos.txt",net0.n_2_2_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_1_yneg.txt",net0.n_2_2_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_1_zpos.txt",net0.n_2_2_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_1_zneg.txt",net0.n_2_2_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_1_xpos.txt",net0.n_2_2_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_1_xneg.txt",net0.n_2_2_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_1_ypos.txt",net0.n_2_2_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_1_yneg.txt",net0.n_2_2_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_1_zpos.txt",net0.n_2_2_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_1_zneg.txt",net0.n_2_2_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_2_local.txt",net0.n_2_2_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_2_xpos.txt",net0.n_2_2_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_2_xneg.txt",net0.n_2_2_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_2_ypos.txt",net0.n_2_2_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_2_yneg.txt",net0.n_2_2_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_2_zpos.txt",net0.n_2_2_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_2_zneg.txt",net0.n_2_2_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_2_xpos.txt",net0.n_2_2_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_2_xneg.txt",net0.n_2_2_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_2_ypos.txt",net0.n_2_2_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_2_yneg.txt",net0.n_2_2_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_2_zpos.txt",net0.n_2_2_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_2_zneg.txt",net0.n_2_2_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_2_xpos.txt",net0.n_2_2_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_2_xneg.txt",net0.n_2_2_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_2_ypos.txt",net0.n_2_2_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_2_yneg.txt",net0.n_2_2_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_2_zpos.txt",net0.n_2_2_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_2_zneg.txt",net0.n_2_2_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_3_local.txt",net0.n_2_2_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_3_xpos.txt",net0.n_2_2_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_3_xneg.txt",net0.n_2_2_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_3_ypos.txt",net0.n_2_2_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_3_yneg.txt",net0.n_2_2_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_3_zpos.txt",net0.n_2_2_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_3_zneg.txt",net0.n_2_2_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_3_xpos.txt",net0.n_2_2_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_3_xneg.txt",net0.n_2_2_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_3_ypos.txt",net0.n_2_2_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_3_yneg.txt",net0.n_2_2_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_3_zpos.txt",net0.n_2_2_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_3_zneg.txt",net0.n_2_2_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_3_xpos.txt",net0.n_2_2_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_3_xneg.txt",net0.n_2_2_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_3_ypos.txt",net0.n_2_2_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_3_yneg.txt",net0.n_2_2_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_3_zpos.txt",net0.n_2_2_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_3_zneg.txt",net0.n_2_2_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_4_local.txt",net0.n_2_2_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_4_xpos.txt",net0.n_2_2_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_4_xneg.txt",net0.n_2_2_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_4_ypos.txt",net0.n_2_2_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_4_yneg.txt",net0.n_2_2_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_4_zpos.txt",net0.n_2_2_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_4_zneg.txt",net0.n_2_2_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_4_xpos.txt",net0.n_2_2_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_4_xneg.txt",net0.n_2_2_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_4_ypos.txt",net0.n_2_2_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_4_yneg.txt",net0.n_2_2_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_4_zpos.txt",net0.n_2_2_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_4_zneg.txt",net0.n_2_2_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_4_xpos.txt",net0.n_2_2_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_4_xneg.txt",net0.n_2_2_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_4_ypos.txt",net0.n_2_2_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_4_yneg.txt",net0.n_2_2_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_4_zpos.txt",net0.n_2_2_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_4_zneg.txt",net0.n_2_2_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_5_local.txt",net0.n_2_2_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_5_xpos.txt",net0.n_2_2_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_5_xneg.txt",net0.n_2_2_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_5_ypos.txt",net0.n_2_2_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_5_yneg.txt",net0.n_2_2_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_5_zpos.txt",net0.n_2_2_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_5_zneg.txt",net0.n_2_2_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_5_xpos.txt",net0.n_2_2_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_5_xneg.txt",net0.n_2_2_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_5_ypos.txt",net0.n_2_2_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_5_yneg.txt",net0.n_2_2_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_5_zpos.txt",net0.n_2_2_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_5_zneg.txt",net0.n_2_2_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_5_xpos.txt",net0.n_2_2_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_5_xneg.txt",net0.n_2_2_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_5_ypos.txt",net0.n_2_2_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_5_yneg.txt",net0.n_2_2_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_5_zpos.txt",net0.n_2_2_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_5_zneg.txt",net0.n_2_2_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_6_local.txt",net0.n_2_2_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_6_xpos.txt",net0.n_2_2_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_6_xneg.txt",net0.n_2_2_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_6_ypos.txt",net0.n_2_2_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_6_yneg.txt",net0.n_2_2_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_6_zpos.txt",net0.n_2_2_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_6_zneg.txt",net0.n_2_2_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_6_xpos.txt",net0.n_2_2_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_6_xneg.txt",net0.n_2_2_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_6_ypos.txt",net0.n_2_2_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_6_yneg.txt",net0.n_2_2_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_6_zpos.txt",net0.n_2_2_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_6_zneg.txt",net0.n_2_2_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_6_xpos.txt",net0.n_2_2_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_6_xneg.txt",net0.n_2_2_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_6_ypos.txt",net0.n_2_2_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_6_yneg.txt",net0.n_2_2_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_6_zpos.txt",net0.n_2_2_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_6_zneg.txt",net0.n_2_2_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_7_local.txt",net0.n_2_2_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_7_xpos.txt",net0.n_2_2_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_7_xneg.txt",net0.n_2_2_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_7_ypos.txt",net0.n_2_2_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_7_yneg.txt",net0.n_2_2_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_7_zpos.txt",net0.n_2_2_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_2_7_zneg.txt",net0.n_2_2_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_7_xpos.txt",net0.n_2_2_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_7_xneg.txt",net0.n_2_2_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_7_ypos.txt",net0.n_2_2_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_7_yneg.txt",net0.n_2_2_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_7_zpos.txt",net0.n_2_2_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_2_7_zneg.txt",net0.n_2_2_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_7_xpos.txt",net0.n_2_2_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_7_xneg.txt",net0.n_2_2_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_7_ypos.txt",net0.n_2_2_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_7_yneg.txt",net0.n_2_2_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_7_zpos.txt",net0.n_2_2_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_2_7_zneg.txt",net0.n_2_2_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_0_local.txt",net0.n_2_3_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_0_xpos.txt",net0.n_2_3_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_0_xneg.txt",net0.n_2_3_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_0_ypos.txt",net0.n_2_3_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_0_yneg.txt",net0.n_2_3_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_0_zpos.txt",net0.n_2_3_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_0_zneg.txt",net0.n_2_3_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_0_xpos.txt",net0.n_2_3_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_0_xneg.txt",net0.n_2_3_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_0_ypos.txt",net0.n_2_3_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_0_yneg.txt",net0.n_2_3_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_0_zpos.txt",net0.n_2_3_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_0_zneg.txt",net0.n_2_3_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_0_xpos.txt",net0.n_2_3_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_0_xneg.txt",net0.n_2_3_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_0_ypos.txt",net0.n_2_3_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_0_yneg.txt",net0.n_2_3_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_0_zpos.txt",net0.n_2_3_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_0_zneg.txt",net0.n_2_3_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_1_local.txt",net0.n_2_3_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_1_xpos.txt",net0.n_2_3_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_1_xneg.txt",net0.n_2_3_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_1_ypos.txt",net0.n_2_3_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_1_yneg.txt",net0.n_2_3_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_1_zpos.txt",net0.n_2_3_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_1_zneg.txt",net0.n_2_3_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_1_xpos.txt",net0.n_2_3_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_1_xneg.txt",net0.n_2_3_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_1_ypos.txt",net0.n_2_3_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_1_yneg.txt",net0.n_2_3_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_1_zpos.txt",net0.n_2_3_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_1_zneg.txt",net0.n_2_3_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_1_xpos.txt",net0.n_2_3_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_1_xneg.txt",net0.n_2_3_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_1_ypos.txt",net0.n_2_3_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_1_yneg.txt",net0.n_2_3_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_1_zpos.txt",net0.n_2_3_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_1_zneg.txt",net0.n_2_3_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_2_local.txt",net0.n_2_3_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_2_xpos.txt",net0.n_2_3_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_2_xneg.txt",net0.n_2_3_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_2_ypos.txt",net0.n_2_3_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_2_yneg.txt",net0.n_2_3_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_2_zpos.txt",net0.n_2_3_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_2_zneg.txt",net0.n_2_3_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_2_xpos.txt",net0.n_2_3_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_2_xneg.txt",net0.n_2_3_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_2_ypos.txt",net0.n_2_3_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_2_yneg.txt",net0.n_2_3_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_2_zpos.txt",net0.n_2_3_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_2_zneg.txt",net0.n_2_3_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_2_xpos.txt",net0.n_2_3_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_2_xneg.txt",net0.n_2_3_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_2_ypos.txt",net0.n_2_3_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_2_yneg.txt",net0.n_2_3_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_2_zpos.txt",net0.n_2_3_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_2_zneg.txt",net0.n_2_3_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_3_local.txt",net0.n_2_3_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_3_xpos.txt",net0.n_2_3_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_3_xneg.txt",net0.n_2_3_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_3_ypos.txt",net0.n_2_3_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_3_yneg.txt",net0.n_2_3_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_3_zpos.txt",net0.n_2_3_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_3_zneg.txt",net0.n_2_3_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_3_xpos.txt",net0.n_2_3_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_3_xneg.txt",net0.n_2_3_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_3_ypos.txt",net0.n_2_3_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_3_yneg.txt",net0.n_2_3_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_3_zpos.txt",net0.n_2_3_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_3_zneg.txt",net0.n_2_3_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_3_xpos.txt",net0.n_2_3_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_3_xneg.txt",net0.n_2_3_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_3_ypos.txt",net0.n_2_3_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_3_yneg.txt",net0.n_2_3_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_3_zpos.txt",net0.n_2_3_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_3_zneg.txt",net0.n_2_3_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_4_local.txt",net0.n_2_3_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_4_xpos.txt",net0.n_2_3_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_4_xneg.txt",net0.n_2_3_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_4_ypos.txt",net0.n_2_3_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_4_yneg.txt",net0.n_2_3_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_4_zpos.txt",net0.n_2_3_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_4_zneg.txt",net0.n_2_3_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_4_xpos.txt",net0.n_2_3_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_4_xneg.txt",net0.n_2_3_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_4_ypos.txt",net0.n_2_3_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_4_yneg.txt",net0.n_2_3_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_4_zpos.txt",net0.n_2_3_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_4_zneg.txt",net0.n_2_3_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_4_xpos.txt",net0.n_2_3_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_4_xneg.txt",net0.n_2_3_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_4_ypos.txt",net0.n_2_3_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_4_yneg.txt",net0.n_2_3_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_4_zpos.txt",net0.n_2_3_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_4_zneg.txt",net0.n_2_3_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_5_local.txt",net0.n_2_3_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_5_xpos.txt",net0.n_2_3_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_5_xneg.txt",net0.n_2_3_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_5_ypos.txt",net0.n_2_3_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_5_yneg.txt",net0.n_2_3_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_5_zpos.txt",net0.n_2_3_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_5_zneg.txt",net0.n_2_3_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_5_xpos.txt",net0.n_2_3_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_5_xneg.txt",net0.n_2_3_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_5_ypos.txt",net0.n_2_3_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_5_yneg.txt",net0.n_2_3_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_5_zpos.txt",net0.n_2_3_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_5_zneg.txt",net0.n_2_3_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_5_xpos.txt",net0.n_2_3_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_5_xneg.txt",net0.n_2_3_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_5_ypos.txt",net0.n_2_3_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_5_yneg.txt",net0.n_2_3_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_5_zpos.txt",net0.n_2_3_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_5_zneg.txt",net0.n_2_3_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_6_local.txt",net0.n_2_3_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_6_xpos.txt",net0.n_2_3_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_6_xneg.txt",net0.n_2_3_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_6_ypos.txt",net0.n_2_3_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_6_yneg.txt",net0.n_2_3_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_6_zpos.txt",net0.n_2_3_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_6_zneg.txt",net0.n_2_3_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_6_xpos.txt",net0.n_2_3_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_6_xneg.txt",net0.n_2_3_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_6_ypos.txt",net0.n_2_3_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_6_yneg.txt",net0.n_2_3_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_6_zpos.txt",net0.n_2_3_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_6_zneg.txt",net0.n_2_3_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_6_xpos.txt",net0.n_2_3_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_6_xneg.txt",net0.n_2_3_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_6_ypos.txt",net0.n_2_3_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_6_yneg.txt",net0.n_2_3_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_6_zpos.txt",net0.n_2_3_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_6_zneg.txt",net0.n_2_3_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_7_local.txt",net0.n_2_3_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_7_xpos.txt",net0.n_2_3_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_7_xneg.txt",net0.n_2_3_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_7_ypos.txt",net0.n_2_3_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_7_yneg.txt",net0.n_2_3_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_7_zpos.txt",net0.n_2_3_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_3_7_zneg.txt",net0.n_2_3_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_7_xpos.txt",net0.n_2_3_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_7_xneg.txt",net0.n_2_3_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_7_ypos.txt",net0.n_2_3_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_7_yneg.txt",net0.n_2_3_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_7_zpos.txt",net0.n_2_3_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_3_7_zneg.txt",net0.n_2_3_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_7_xpos.txt",net0.n_2_3_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_7_xneg.txt",net0.n_2_3_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_7_ypos.txt",net0.n_2_3_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_7_yneg.txt",net0.n_2_3_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_7_zpos.txt",net0.n_2_3_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_3_7_zneg.txt",net0.n_2_3_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_0_local.txt",net0.n_2_4_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_0_xpos.txt",net0.n_2_4_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_0_xneg.txt",net0.n_2_4_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_0_ypos.txt",net0.n_2_4_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_0_yneg.txt",net0.n_2_4_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_0_zpos.txt",net0.n_2_4_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_0_zneg.txt",net0.n_2_4_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_0_xpos.txt",net0.n_2_4_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_0_xneg.txt",net0.n_2_4_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_0_ypos.txt",net0.n_2_4_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_0_yneg.txt",net0.n_2_4_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_0_zpos.txt",net0.n_2_4_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_0_zneg.txt",net0.n_2_4_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_0_xpos.txt",net0.n_2_4_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_0_xneg.txt",net0.n_2_4_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_0_ypos.txt",net0.n_2_4_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_0_yneg.txt",net0.n_2_4_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_0_zpos.txt",net0.n_2_4_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_0_zneg.txt",net0.n_2_4_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_1_local.txt",net0.n_2_4_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_1_xpos.txt",net0.n_2_4_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_1_xneg.txt",net0.n_2_4_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_1_ypos.txt",net0.n_2_4_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_1_yneg.txt",net0.n_2_4_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_1_zpos.txt",net0.n_2_4_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_1_zneg.txt",net0.n_2_4_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_1_xpos.txt",net0.n_2_4_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_1_xneg.txt",net0.n_2_4_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_1_ypos.txt",net0.n_2_4_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_1_yneg.txt",net0.n_2_4_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_1_zpos.txt",net0.n_2_4_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_1_zneg.txt",net0.n_2_4_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_1_xpos.txt",net0.n_2_4_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_1_xneg.txt",net0.n_2_4_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_1_ypos.txt",net0.n_2_4_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_1_yneg.txt",net0.n_2_4_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_1_zpos.txt",net0.n_2_4_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_1_zneg.txt",net0.n_2_4_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_2_local.txt",net0.n_2_4_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_2_xpos.txt",net0.n_2_4_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_2_xneg.txt",net0.n_2_4_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_2_ypos.txt",net0.n_2_4_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_2_yneg.txt",net0.n_2_4_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_2_zpos.txt",net0.n_2_4_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_2_zneg.txt",net0.n_2_4_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_2_xpos.txt",net0.n_2_4_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_2_xneg.txt",net0.n_2_4_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_2_ypos.txt",net0.n_2_4_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_2_yneg.txt",net0.n_2_4_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_2_zpos.txt",net0.n_2_4_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_2_zneg.txt",net0.n_2_4_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_2_xpos.txt",net0.n_2_4_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_2_xneg.txt",net0.n_2_4_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_2_ypos.txt",net0.n_2_4_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_2_yneg.txt",net0.n_2_4_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_2_zpos.txt",net0.n_2_4_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_2_zneg.txt",net0.n_2_4_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_3_local.txt",net0.n_2_4_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_3_xpos.txt",net0.n_2_4_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_3_xneg.txt",net0.n_2_4_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_3_ypos.txt",net0.n_2_4_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_3_yneg.txt",net0.n_2_4_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_3_zpos.txt",net0.n_2_4_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_3_zneg.txt",net0.n_2_4_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_3_xpos.txt",net0.n_2_4_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_3_xneg.txt",net0.n_2_4_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_3_ypos.txt",net0.n_2_4_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_3_yneg.txt",net0.n_2_4_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_3_zpos.txt",net0.n_2_4_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_3_zneg.txt",net0.n_2_4_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_3_xpos.txt",net0.n_2_4_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_3_xneg.txt",net0.n_2_4_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_3_ypos.txt",net0.n_2_4_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_3_yneg.txt",net0.n_2_4_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_3_zpos.txt",net0.n_2_4_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_3_zneg.txt",net0.n_2_4_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_4_local.txt",net0.n_2_4_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_4_xpos.txt",net0.n_2_4_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_4_xneg.txt",net0.n_2_4_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_4_ypos.txt",net0.n_2_4_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_4_yneg.txt",net0.n_2_4_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_4_zpos.txt",net0.n_2_4_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_4_zneg.txt",net0.n_2_4_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_4_xpos.txt",net0.n_2_4_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_4_xneg.txt",net0.n_2_4_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_4_ypos.txt",net0.n_2_4_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_4_yneg.txt",net0.n_2_4_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_4_zpos.txt",net0.n_2_4_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_4_zneg.txt",net0.n_2_4_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_4_xpos.txt",net0.n_2_4_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_4_xneg.txt",net0.n_2_4_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_4_ypos.txt",net0.n_2_4_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_4_yneg.txt",net0.n_2_4_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_4_zpos.txt",net0.n_2_4_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_4_zneg.txt",net0.n_2_4_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_5_local.txt",net0.n_2_4_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_5_xpos.txt",net0.n_2_4_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_5_xneg.txt",net0.n_2_4_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_5_ypos.txt",net0.n_2_4_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_5_yneg.txt",net0.n_2_4_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_5_zpos.txt",net0.n_2_4_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_5_zneg.txt",net0.n_2_4_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_5_xpos.txt",net0.n_2_4_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_5_xneg.txt",net0.n_2_4_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_5_ypos.txt",net0.n_2_4_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_5_yneg.txt",net0.n_2_4_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_5_zpos.txt",net0.n_2_4_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_5_zneg.txt",net0.n_2_4_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_5_xpos.txt",net0.n_2_4_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_5_xneg.txt",net0.n_2_4_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_5_ypos.txt",net0.n_2_4_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_5_yneg.txt",net0.n_2_4_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_5_zpos.txt",net0.n_2_4_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_5_zneg.txt",net0.n_2_4_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_6_local.txt",net0.n_2_4_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_6_xpos.txt",net0.n_2_4_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_6_xneg.txt",net0.n_2_4_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_6_ypos.txt",net0.n_2_4_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_6_yneg.txt",net0.n_2_4_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_6_zpos.txt",net0.n_2_4_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_6_zneg.txt",net0.n_2_4_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_6_xpos.txt",net0.n_2_4_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_6_xneg.txt",net0.n_2_4_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_6_ypos.txt",net0.n_2_4_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_6_yneg.txt",net0.n_2_4_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_6_zpos.txt",net0.n_2_4_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_6_zneg.txt",net0.n_2_4_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_6_xpos.txt",net0.n_2_4_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_6_xneg.txt",net0.n_2_4_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_6_ypos.txt",net0.n_2_4_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_6_yneg.txt",net0.n_2_4_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_6_zpos.txt",net0.n_2_4_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_6_zneg.txt",net0.n_2_4_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_7_local.txt",net0.n_2_4_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_7_xpos.txt",net0.n_2_4_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_7_xneg.txt",net0.n_2_4_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_7_ypos.txt",net0.n_2_4_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_7_yneg.txt",net0.n_2_4_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_7_zpos.txt",net0.n_2_4_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_4_7_zneg.txt",net0.n_2_4_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_7_xpos.txt",net0.n_2_4_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_7_xneg.txt",net0.n_2_4_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_7_ypos.txt",net0.n_2_4_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_7_yneg.txt",net0.n_2_4_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_7_zpos.txt",net0.n_2_4_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_4_7_zneg.txt",net0.n_2_4_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_7_xpos.txt",net0.n_2_4_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_7_xneg.txt",net0.n_2_4_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_7_ypos.txt",net0.n_2_4_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_7_yneg.txt",net0.n_2_4_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_7_zpos.txt",net0.n_2_4_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_4_7_zneg.txt",net0.n_2_4_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_0_local.txt",net0.n_2_5_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_0_xpos.txt",net0.n_2_5_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_0_xneg.txt",net0.n_2_5_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_0_ypos.txt",net0.n_2_5_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_0_yneg.txt",net0.n_2_5_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_0_zpos.txt",net0.n_2_5_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_0_zneg.txt",net0.n_2_5_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_0_xpos.txt",net0.n_2_5_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_0_xneg.txt",net0.n_2_5_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_0_ypos.txt",net0.n_2_5_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_0_yneg.txt",net0.n_2_5_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_0_zpos.txt",net0.n_2_5_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_0_zneg.txt",net0.n_2_5_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_0_xpos.txt",net0.n_2_5_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_0_xneg.txt",net0.n_2_5_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_0_ypos.txt",net0.n_2_5_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_0_yneg.txt",net0.n_2_5_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_0_zpos.txt",net0.n_2_5_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_0_zneg.txt",net0.n_2_5_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_1_local.txt",net0.n_2_5_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_1_xpos.txt",net0.n_2_5_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_1_xneg.txt",net0.n_2_5_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_1_ypos.txt",net0.n_2_5_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_1_yneg.txt",net0.n_2_5_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_1_zpos.txt",net0.n_2_5_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_1_zneg.txt",net0.n_2_5_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_1_xpos.txt",net0.n_2_5_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_1_xneg.txt",net0.n_2_5_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_1_ypos.txt",net0.n_2_5_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_1_yneg.txt",net0.n_2_5_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_1_zpos.txt",net0.n_2_5_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_1_zneg.txt",net0.n_2_5_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_1_xpos.txt",net0.n_2_5_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_1_xneg.txt",net0.n_2_5_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_1_ypos.txt",net0.n_2_5_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_1_yneg.txt",net0.n_2_5_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_1_zpos.txt",net0.n_2_5_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_1_zneg.txt",net0.n_2_5_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_2_local.txt",net0.n_2_5_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_2_xpos.txt",net0.n_2_5_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_2_xneg.txt",net0.n_2_5_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_2_ypos.txt",net0.n_2_5_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_2_yneg.txt",net0.n_2_5_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_2_zpos.txt",net0.n_2_5_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_2_zneg.txt",net0.n_2_5_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_2_xpos.txt",net0.n_2_5_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_2_xneg.txt",net0.n_2_5_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_2_ypos.txt",net0.n_2_5_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_2_yneg.txt",net0.n_2_5_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_2_zpos.txt",net0.n_2_5_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_2_zneg.txt",net0.n_2_5_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_2_xpos.txt",net0.n_2_5_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_2_xneg.txt",net0.n_2_5_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_2_ypos.txt",net0.n_2_5_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_2_yneg.txt",net0.n_2_5_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_2_zpos.txt",net0.n_2_5_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_2_zneg.txt",net0.n_2_5_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_3_local.txt",net0.n_2_5_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_3_xpos.txt",net0.n_2_5_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_3_xneg.txt",net0.n_2_5_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_3_ypos.txt",net0.n_2_5_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_3_yneg.txt",net0.n_2_5_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_3_zpos.txt",net0.n_2_5_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_3_zneg.txt",net0.n_2_5_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_3_xpos.txt",net0.n_2_5_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_3_xneg.txt",net0.n_2_5_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_3_ypos.txt",net0.n_2_5_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_3_yneg.txt",net0.n_2_5_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_3_zpos.txt",net0.n_2_5_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_3_zneg.txt",net0.n_2_5_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_3_xpos.txt",net0.n_2_5_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_3_xneg.txt",net0.n_2_5_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_3_ypos.txt",net0.n_2_5_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_3_yneg.txt",net0.n_2_5_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_3_zpos.txt",net0.n_2_5_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_3_zneg.txt",net0.n_2_5_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_4_local.txt",net0.n_2_5_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_4_xpos.txt",net0.n_2_5_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_4_xneg.txt",net0.n_2_5_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_4_ypos.txt",net0.n_2_5_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_4_yneg.txt",net0.n_2_5_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_4_zpos.txt",net0.n_2_5_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_4_zneg.txt",net0.n_2_5_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_4_xpos.txt",net0.n_2_5_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_4_xneg.txt",net0.n_2_5_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_4_ypos.txt",net0.n_2_5_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_4_yneg.txt",net0.n_2_5_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_4_zpos.txt",net0.n_2_5_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_4_zneg.txt",net0.n_2_5_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_4_xpos.txt",net0.n_2_5_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_4_xneg.txt",net0.n_2_5_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_4_ypos.txt",net0.n_2_5_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_4_yneg.txt",net0.n_2_5_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_4_zpos.txt",net0.n_2_5_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_4_zneg.txt",net0.n_2_5_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_5_local.txt",net0.n_2_5_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_5_xpos.txt",net0.n_2_5_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_5_xneg.txt",net0.n_2_5_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_5_ypos.txt",net0.n_2_5_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_5_yneg.txt",net0.n_2_5_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_5_zpos.txt",net0.n_2_5_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_5_zneg.txt",net0.n_2_5_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_5_xpos.txt",net0.n_2_5_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_5_xneg.txt",net0.n_2_5_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_5_ypos.txt",net0.n_2_5_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_5_yneg.txt",net0.n_2_5_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_5_zpos.txt",net0.n_2_5_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_5_zneg.txt",net0.n_2_5_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_5_xpos.txt",net0.n_2_5_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_5_xneg.txt",net0.n_2_5_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_5_ypos.txt",net0.n_2_5_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_5_yneg.txt",net0.n_2_5_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_5_zpos.txt",net0.n_2_5_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_5_zneg.txt",net0.n_2_5_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_6_local.txt",net0.n_2_5_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_6_xpos.txt",net0.n_2_5_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_6_xneg.txt",net0.n_2_5_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_6_ypos.txt",net0.n_2_5_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_6_yneg.txt",net0.n_2_5_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_6_zpos.txt",net0.n_2_5_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_6_zneg.txt",net0.n_2_5_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_6_xpos.txt",net0.n_2_5_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_6_xneg.txt",net0.n_2_5_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_6_ypos.txt",net0.n_2_5_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_6_yneg.txt",net0.n_2_5_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_6_zpos.txt",net0.n_2_5_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_6_zneg.txt",net0.n_2_5_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_6_xpos.txt",net0.n_2_5_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_6_xneg.txt",net0.n_2_5_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_6_ypos.txt",net0.n_2_5_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_6_yneg.txt",net0.n_2_5_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_6_zpos.txt",net0.n_2_5_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_6_zneg.txt",net0.n_2_5_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_7_local.txt",net0.n_2_5_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_7_xpos.txt",net0.n_2_5_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_7_xneg.txt",net0.n_2_5_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_7_ypos.txt",net0.n_2_5_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_7_yneg.txt",net0.n_2_5_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_7_zpos.txt",net0.n_2_5_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_5_7_zneg.txt",net0.n_2_5_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_7_xpos.txt",net0.n_2_5_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_7_xneg.txt",net0.n_2_5_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_7_ypos.txt",net0.n_2_5_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_7_yneg.txt",net0.n_2_5_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_7_zpos.txt",net0.n_2_5_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_5_7_zneg.txt",net0.n_2_5_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_7_xpos.txt",net0.n_2_5_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_7_xneg.txt",net0.n_2_5_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_7_ypos.txt",net0.n_2_5_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_7_yneg.txt",net0.n_2_5_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_7_zpos.txt",net0.n_2_5_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_5_7_zneg.txt",net0.n_2_5_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_0_local.txt",net0.n_2_6_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_0_xpos.txt",net0.n_2_6_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_0_xneg.txt",net0.n_2_6_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_0_ypos.txt",net0.n_2_6_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_0_yneg.txt",net0.n_2_6_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_0_zpos.txt",net0.n_2_6_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_0_zneg.txt",net0.n_2_6_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_0_xpos.txt",net0.n_2_6_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_0_xneg.txt",net0.n_2_6_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_0_ypos.txt",net0.n_2_6_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_0_yneg.txt",net0.n_2_6_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_0_zpos.txt",net0.n_2_6_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_0_zneg.txt",net0.n_2_6_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_0_xpos.txt",net0.n_2_6_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_0_xneg.txt",net0.n_2_6_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_0_ypos.txt",net0.n_2_6_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_0_yneg.txt",net0.n_2_6_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_0_zpos.txt",net0.n_2_6_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_0_zneg.txt",net0.n_2_6_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_1_local.txt",net0.n_2_6_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_1_xpos.txt",net0.n_2_6_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_1_xneg.txt",net0.n_2_6_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_1_ypos.txt",net0.n_2_6_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_1_yneg.txt",net0.n_2_6_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_1_zpos.txt",net0.n_2_6_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_1_zneg.txt",net0.n_2_6_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_1_xpos.txt",net0.n_2_6_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_1_xneg.txt",net0.n_2_6_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_1_ypos.txt",net0.n_2_6_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_1_yneg.txt",net0.n_2_6_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_1_zpos.txt",net0.n_2_6_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_1_zneg.txt",net0.n_2_6_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_1_xpos.txt",net0.n_2_6_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_1_xneg.txt",net0.n_2_6_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_1_ypos.txt",net0.n_2_6_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_1_yneg.txt",net0.n_2_6_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_1_zpos.txt",net0.n_2_6_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_1_zneg.txt",net0.n_2_6_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_2_local.txt",net0.n_2_6_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_2_xpos.txt",net0.n_2_6_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_2_xneg.txt",net0.n_2_6_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_2_ypos.txt",net0.n_2_6_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_2_yneg.txt",net0.n_2_6_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_2_zpos.txt",net0.n_2_6_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_2_zneg.txt",net0.n_2_6_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_2_xpos.txt",net0.n_2_6_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_2_xneg.txt",net0.n_2_6_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_2_ypos.txt",net0.n_2_6_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_2_yneg.txt",net0.n_2_6_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_2_zpos.txt",net0.n_2_6_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_2_zneg.txt",net0.n_2_6_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_2_xpos.txt",net0.n_2_6_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_2_xneg.txt",net0.n_2_6_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_2_ypos.txt",net0.n_2_6_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_2_yneg.txt",net0.n_2_6_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_2_zpos.txt",net0.n_2_6_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_2_zneg.txt",net0.n_2_6_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_3_local.txt",net0.n_2_6_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_3_xpos.txt",net0.n_2_6_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_3_xneg.txt",net0.n_2_6_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_3_ypos.txt",net0.n_2_6_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_3_yneg.txt",net0.n_2_6_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_3_zpos.txt",net0.n_2_6_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_3_zneg.txt",net0.n_2_6_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_3_xpos.txt",net0.n_2_6_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_3_xneg.txt",net0.n_2_6_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_3_ypos.txt",net0.n_2_6_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_3_yneg.txt",net0.n_2_6_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_3_zpos.txt",net0.n_2_6_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_3_zneg.txt",net0.n_2_6_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_3_xpos.txt",net0.n_2_6_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_3_xneg.txt",net0.n_2_6_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_3_ypos.txt",net0.n_2_6_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_3_yneg.txt",net0.n_2_6_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_3_zpos.txt",net0.n_2_6_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_3_zneg.txt",net0.n_2_6_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_4_local.txt",net0.n_2_6_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_4_xpos.txt",net0.n_2_6_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_4_xneg.txt",net0.n_2_6_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_4_ypos.txt",net0.n_2_6_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_4_yneg.txt",net0.n_2_6_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_4_zpos.txt",net0.n_2_6_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_4_zneg.txt",net0.n_2_6_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_4_xpos.txt",net0.n_2_6_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_4_xneg.txt",net0.n_2_6_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_4_ypos.txt",net0.n_2_6_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_4_yneg.txt",net0.n_2_6_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_4_zpos.txt",net0.n_2_6_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_4_zneg.txt",net0.n_2_6_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_4_xpos.txt",net0.n_2_6_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_4_xneg.txt",net0.n_2_6_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_4_ypos.txt",net0.n_2_6_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_4_yneg.txt",net0.n_2_6_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_4_zpos.txt",net0.n_2_6_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_4_zneg.txt",net0.n_2_6_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_5_local.txt",net0.n_2_6_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_5_xpos.txt",net0.n_2_6_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_5_xneg.txt",net0.n_2_6_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_5_ypos.txt",net0.n_2_6_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_5_yneg.txt",net0.n_2_6_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_5_zpos.txt",net0.n_2_6_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_5_zneg.txt",net0.n_2_6_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_5_xpos.txt",net0.n_2_6_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_5_xneg.txt",net0.n_2_6_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_5_ypos.txt",net0.n_2_6_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_5_yneg.txt",net0.n_2_6_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_5_zpos.txt",net0.n_2_6_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_5_zneg.txt",net0.n_2_6_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_5_xpos.txt",net0.n_2_6_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_5_xneg.txt",net0.n_2_6_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_5_ypos.txt",net0.n_2_6_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_5_yneg.txt",net0.n_2_6_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_5_zpos.txt",net0.n_2_6_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_5_zneg.txt",net0.n_2_6_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_6_local.txt",net0.n_2_6_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_6_xpos.txt",net0.n_2_6_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_6_xneg.txt",net0.n_2_6_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_6_ypos.txt",net0.n_2_6_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_6_yneg.txt",net0.n_2_6_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_6_zpos.txt",net0.n_2_6_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_6_zneg.txt",net0.n_2_6_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_6_xpos.txt",net0.n_2_6_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_6_xneg.txt",net0.n_2_6_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_6_ypos.txt",net0.n_2_6_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_6_yneg.txt",net0.n_2_6_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_6_zpos.txt",net0.n_2_6_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_6_zneg.txt",net0.n_2_6_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_6_xpos.txt",net0.n_2_6_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_6_xneg.txt",net0.n_2_6_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_6_ypos.txt",net0.n_2_6_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_6_yneg.txt",net0.n_2_6_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_6_zpos.txt",net0.n_2_6_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_6_zneg.txt",net0.n_2_6_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_7_local.txt",net0.n_2_6_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_7_xpos.txt",net0.n_2_6_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_7_xneg.txt",net0.n_2_6_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_7_ypos.txt",net0.n_2_6_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_7_yneg.txt",net0.n_2_6_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_7_zpos.txt",net0.n_2_6_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_6_7_zneg.txt",net0.n_2_6_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_7_xpos.txt",net0.n_2_6_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_7_xneg.txt",net0.n_2_6_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_7_ypos.txt",net0.n_2_6_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_7_yneg.txt",net0.n_2_6_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_7_zpos.txt",net0.n_2_6_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_6_7_zneg.txt",net0.n_2_6_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_7_xpos.txt",net0.n_2_6_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_7_xneg.txt",net0.n_2_6_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_7_ypos.txt",net0.n_2_6_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_7_yneg.txt",net0.n_2_6_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_7_zpos.txt",net0.n_2_6_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_6_7_zneg.txt",net0.n_2_6_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_0_local.txt",net0.n_2_7_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_0_xpos.txt",net0.n_2_7_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_0_xneg.txt",net0.n_2_7_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_0_ypos.txt",net0.n_2_7_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_0_yneg.txt",net0.n_2_7_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_0_zpos.txt",net0.n_2_7_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_0_zneg.txt",net0.n_2_7_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_0_xpos.txt",net0.n_2_7_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_0_xneg.txt",net0.n_2_7_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_0_ypos.txt",net0.n_2_7_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_0_yneg.txt",net0.n_2_7_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_0_zpos.txt",net0.n_2_7_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_0_zneg.txt",net0.n_2_7_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_0_xpos.txt",net0.n_2_7_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_0_xneg.txt",net0.n_2_7_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_0_ypos.txt",net0.n_2_7_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_0_yneg.txt",net0.n_2_7_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_0_zpos.txt",net0.n_2_7_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_0_zneg.txt",net0.n_2_7_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_1_local.txt",net0.n_2_7_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_1_xpos.txt",net0.n_2_7_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_1_xneg.txt",net0.n_2_7_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_1_ypos.txt",net0.n_2_7_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_1_yneg.txt",net0.n_2_7_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_1_zpos.txt",net0.n_2_7_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_1_zneg.txt",net0.n_2_7_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_1_xpos.txt",net0.n_2_7_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_1_xneg.txt",net0.n_2_7_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_1_ypos.txt",net0.n_2_7_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_1_yneg.txt",net0.n_2_7_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_1_zpos.txt",net0.n_2_7_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_1_zneg.txt",net0.n_2_7_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_1_xpos.txt",net0.n_2_7_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_1_xneg.txt",net0.n_2_7_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_1_ypos.txt",net0.n_2_7_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_1_yneg.txt",net0.n_2_7_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_1_zpos.txt",net0.n_2_7_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_1_zneg.txt",net0.n_2_7_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_2_local.txt",net0.n_2_7_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_2_xpos.txt",net0.n_2_7_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_2_xneg.txt",net0.n_2_7_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_2_ypos.txt",net0.n_2_7_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_2_yneg.txt",net0.n_2_7_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_2_zpos.txt",net0.n_2_7_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_2_zneg.txt",net0.n_2_7_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_2_xpos.txt",net0.n_2_7_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_2_xneg.txt",net0.n_2_7_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_2_ypos.txt",net0.n_2_7_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_2_yneg.txt",net0.n_2_7_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_2_zpos.txt",net0.n_2_7_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_2_zneg.txt",net0.n_2_7_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_2_xpos.txt",net0.n_2_7_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_2_xneg.txt",net0.n_2_7_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_2_ypos.txt",net0.n_2_7_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_2_yneg.txt",net0.n_2_7_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_2_zpos.txt",net0.n_2_7_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_2_zneg.txt",net0.n_2_7_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_3_local.txt",net0.n_2_7_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_3_xpos.txt",net0.n_2_7_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_3_xneg.txt",net0.n_2_7_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_3_ypos.txt",net0.n_2_7_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_3_yneg.txt",net0.n_2_7_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_3_zpos.txt",net0.n_2_7_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_3_zneg.txt",net0.n_2_7_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_3_xpos.txt",net0.n_2_7_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_3_xneg.txt",net0.n_2_7_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_3_ypos.txt",net0.n_2_7_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_3_yneg.txt",net0.n_2_7_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_3_zpos.txt",net0.n_2_7_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_3_zneg.txt",net0.n_2_7_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_3_xpos.txt",net0.n_2_7_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_3_xneg.txt",net0.n_2_7_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_3_ypos.txt",net0.n_2_7_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_3_yneg.txt",net0.n_2_7_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_3_zpos.txt",net0.n_2_7_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_3_zneg.txt",net0.n_2_7_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_4_local.txt",net0.n_2_7_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_4_xpos.txt",net0.n_2_7_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_4_xneg.txt",net0.n_2_7_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_4_ypos.txt",net0.n_2_7_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_4_yneg.txt",net0.n_2_7_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_4_zpos.txt",net0.n_2_7_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_4_zneg.txt",net0.n_2_7_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_4_xpos.txt",net0.n_2_7_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_4_xneg.txt",net0.n_2_7_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_4_ypos.txt",net0.n_2_7_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_4_yneg.txt",net0.n_2_7_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_4_zpos.txt",net0.n_2_7_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_4_zneg.txt",net0.n_2_7_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_4_xpos.txt",net0.n_2_7_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_4_xneg.txt",net0.n_2_7_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_4_ypos.txt",net0.n_2_7_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_4_yneg.txt",net0.n_2_7_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_4_zpos.txt",net0.n_2_7_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_4_zneg.txt",net0.n_2_7_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_5_local.txt",net0.n_2_7_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_5_xpos.txt",net0.n_2_7_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_5_xneg.txt",net0.n_2_7_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_5_ypos.txt",net0.n_2_7_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_5_yneg.txt",net0.n_2_7_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_5_zpos.txt",net0.n_2_7_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_5_zneg.txt",net0.n_2_7_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_5_xpos.txt",net0.n_2_7_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_5_xneg.txt",net0.n_2_7_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_5_ypos.txt",net0.n_2_7_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_5_yneg.txt",net0.n_2_7_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_5_zpos.txt",net0.n_2_7_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_5_zneg.txt",net0.n_2_7_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_5_xpos.txt",net0.n_2_7_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_5_xneg.txt",net0.n_2_7_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_5_ypos.txt",net0.n_2_7_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_5_yneg.txt",net0.n_2_7_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_5_zpos.txt",net0.n_2_7_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_5_zneg.txt",net0.n_2_7_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_6_local.txt",net0.n_2_7_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_6_xpos.txt",net0.n_2_7_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_6_xneg.txt",net0.n_2_7_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_6_ypos.txt",net0.n_2_7_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_6_yneg.txt",net0.n_2_7_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_6_zpos.txt",net0.n_2_7_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_6_zneg.txt",net0.n_2_7_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_6_xpos.txt",net0.n_2_7_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_6_xneg.txt",net0.n_2_7_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_6_ypos.txt",net0.n_2_7_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_6_yneg.txt",net0.n_2_7_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_6_zpos.txt",net0.n_2_7_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_6_zneg.txt",net0.n_2_7_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_6_xpos.txt",net0.n_2_7_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_6_xneg.txt",net0.n_2_7_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_6_ypos.txt",net0.n_2_7_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_6_yneg.txt",net0.n_2_7_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_6_zpos.txt",net0.n_2_7_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_6_zneg.txt",net0.n_2_7_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_7_local.txt",net0.n_2_7_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_7_xpos.txt",net0.n_2_7_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_7_xneg.txt",net0.n_2_7_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_7_ypos.txt",net0.n_2_7_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_7_yneg.txt",net0.n_2_7_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_7_zpos.txt",net0.n_2_7_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_2_7_7_zneg.txt",net0.n_2_7_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_7_xpos.txt",net0.n_2_7_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_7_xneg.txt",net0.n_2_7_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_7_ypos.txt",net0.n_2_7_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_7_yneg.txt",net0.n_2_7_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_7_zpos.txt",net0.n_2_7_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_2_7_7_zneg.txt",net0.n_2_7_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_7_xpos.txt",net0.n_2_7_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_7_xneg.txt",net0.n_2_7_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_7_ypos.txt",net0.n_2_7_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_7_yneg.txt",net0.n_2_7_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_7_zpos.txt",net0.n_2_7_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_2_7_7_zneg.txt",net0.n_2_7_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_0_local.txt",net0.n_3_0_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_0_xpos.txt",net0.n_3_0_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_0_xneg.txt",net0.n_3_0_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_0_ypos.txt",net0.n_3_0_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_0_yneg.txt",net0.n_3_0_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_0_zpos.txt",net0.n_3_0_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_0_zneg.txt",net0.n_3_0_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_0_xpos.txt",net0.n_3_0_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_0_xneg.txt",net0.n_3_0_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_0_ypos.txt",net0.n_3_0_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_0_yneg.txt",net0.n_3_0_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_0_zpos.txt",net0.n_3_0_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_0_zneg.txt",net0.n_3_0_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_0_xpos.txt",net0.n_3_0_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_0_xneg.txt",net0.n_3_0_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_0_ypos.txt",net0.n_3_0_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_0_yneg.txt",net0.n_3_0_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_0_zpos.txt",net0.n_3_0_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_0_zneg.txt",net0.n_3_0_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_1_local.txt",net0.n_3_0_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_1_xpos.txt",net0.n_3_0_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_1_xneg.txt",net0.n_3_0_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_1_ypos.txt",net0.n_3_0_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_1_yneg.txt",net0.n_3_0_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_1_zpos.txt",net0.n_3_0_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_1_zneg.txt",net0.n_3_0_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_1_xpos.txt",net0.n_3_0_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_1_xneg.txt",net0.n_3_0_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_1_ypos.txt",net0.n_3_0_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_1_yneg.txt",net0.n_3_0_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_1_zpos.txt",net0.n_3_0_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_1_zneg.txt",net0.n_3_0_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_1_xpos.txt",net0.n_3_0_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_1_xneg.txt",net0.n_3_0_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_1_ypos.txt",net0.n_3_0_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_1_yneg.txt",net0.n_3_0_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_1_zpos.txt",net0.n_3_0_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_1_zneg.txt",net0.n_3_0_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_2_local.txt",net0.n_3_0_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_2_xpos.txt",net0.n_3_0_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_2_xneg.txt",net0.n_3_0_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_2_ypos.txt",net0.n_3_0_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_2_yneg.txt",net0.n_3_0_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_2_zpos.txt",net0.n_3_0_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_2_zneg.txt",net0.n_3_0_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_2_xpos.txt",net0.n_3_0_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_2_xneg.txt",net0.n_3_0_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_2_ypos.txt",net0.n_3_0_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_2_yneg.txt",net0.n_3_0_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_2_zpos.txt",net0.n_3_0_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_2_zneg.txt",net0.n_3_0_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_2_xpos.txt",net0.n_3_0_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_2_xneg.txt",net0.n_3_0_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_2_ypos.txt",net0.n_3_0_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_2_yneg.txt",net0.n_3_0_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_2_zpos.txt",net0.n_3_0_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_2_zneg.txt",net0.n_3_0_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_3_local.txt",net0.n_3_0_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_3_xpos.txt",net0.n_3_0_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_3_xneg.txt",net0.n_3_0_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_3_ypos.txt",net0.n_3_0_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_3_yneg.txt",net0.n_3_0_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_3_zpos.txt",net0.n_3_0_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_3_zneg.txt",net0.n_3_0_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_3_xpos.txt",net0.n_3_0_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_3_xneg.txt",net0.n_3_0_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_3_ypos.txt",net0.n_3_0_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_3_yneg.txt",net0.n_3_0_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_3_zpos.txt",net0.n_3_0_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_3_zneg.txt",net0.n_3_0_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_3_xpos.txt",net0.n_3_0_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_3_xneg.txt",net0.n_3_0_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_3_ypos.txt",net0.n_3_0_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_3_yneg.txt",net0.n_3_0_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_3_zpos.txt",net0.n_3_0_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_3_zneg.txt",net0.n_3_0_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_4_local.txt",net0.n_3_0_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_4_xpos.txt",net0.n_3_0_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_4_xneg.txt",net0.n_3_0_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_4_ypos.txt",net0.n_3_0_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_4_yneg.txt",net0.n_3_0_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_4_zpos.txt",net0.n_3_0_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_4_zneg.txt",net0.n_3_0_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_4_xpos.txt",net0.n_3_0_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_4_xneg.txt",net0.n_3_0_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_4_ypos.txt",net0.n_3_0_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_4_yneg.txt",net0.n_3_0_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_4_zpos.txt",net0.n_3_0_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_4_zneg.txt",net0.n_3_0_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_4_xpos.txt",net0.n_3_0_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_4_xneg.txt",net0.n_3_0_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_4_ypos.txt",net0.n_3_0_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_4_yneg.txt",net0.n_3_0_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_4_zpos.txt",net0.n_3_0_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_4_zneg.txt",net0.n_3_0_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_5_local.txt",net0.n_3_0_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_5_xpos.txt",net0.n_3_0_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_5_xneg.txt",net0.n_3_0_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_5_ypos.txt",net0.n_3_0_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_5_yneg.txt",net0.n_3_0_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_5_zpos.txt",net0.n_3_0_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_5_zneg.txt",net0.n_3_0_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_5_xpos.txt",net0.n_3_0_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_5_xneg.txt",net0.n_3_0_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_5_ypos.txt",net0.n_3_0_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_5_yneg.txt",net0.n_3_0_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_5_zpos.txt",net0.n_3_0_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_5_zneg.txt",net0.n_3_0_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_5_xpos.txt",net0.n_3_0_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_5_xneg.txt",net0.n_3_0_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_5_ypos.txt",net0.n_3_0_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_5_yneg.txt",net0.n_3_0_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_5_zpos.txt",net0.n_3_0_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_5_zneg.txt",net0.n_3_0_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_6_local.txt",net0.n_3_0_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_6_xpos.txt",net0.n_3_0_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_6_xneg.txt",net0.n_3_0_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_6_ypos.txt",net0.n_3_0_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_6_yneg.txt",net0.n_3_0_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_6_zpos.txt",net0.n_3_0_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_6_zneg.txt",net0.n_3_0_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_6_xpos.txt",net0.n_3_0_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_6_xneg.txt",net0.n_3_0_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_6_ypos.txt",net0.n_3_0_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_6_yneg.txt",net0.n_3_0_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_6_zpos.txt",net0.n_3_0_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_6_zneg.txt",net0.n_3_0_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_6_xpos.txt",net0.n_3_0_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_6_xneg.txt",net0.n_3_0_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_6_ypos.txt",net0.n_3_0_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_6_yneg.txt",net0.n_3_0_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_6_zpos.txt",net0.n_3_0_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_6_zneg.txt",net0.n_3_0_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_7_local.txt",net0.n_3_0_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_7_xpos.txt",net0.n_3_0_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_7_xneg.txt",net0.n_3_0_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_7_ypos.txt",net0.n_3_0_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_7_yneg.txt",net0.n_3_0_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_7_zpos.txt",net0.n_3_0_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_0_7_zneg.txt",net0.n_3_0_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_7_xpos.txt",net0.n_3_0_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_7_xneg.txt",net0.n_3_0_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_7_ypos.txt",net0.n_3_0_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_7_yneg.txt",net0.n_3_0_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_7_zpos.txt",net0.n_3_0_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_0_7_zneg.txt",net0.n_3_0_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_7_xpos.txt",net0.n_3_0_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_7_xneg.txt",net0.n_3_0_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_7_ypos.txt",net0.n_3_0_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_7_yneg.txt",net0.n_3_0_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_7_zpos.txt",net0.n_3_0_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_0_7_zneg.txt",net0.n_3_0_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_0_local.txt",net0.n_3_1_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_0_xpos.txt",net0.n_3_1_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_0_xneg.txt",net0.n_3_1_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_0_ypos.txt",net0.n_3_1_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_0_yneg.txt",net0.n_3_1_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_0_zpos.txt",net0.n_3_1_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_0_zneg.txt",net0.n_3_1_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_0_xpos.txt",net0.n_3_1_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_0_xneg.txt",net0.n_3_1_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_0_ypos.txt",net0.n_3_1_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_0_yneg.txt",net0.n_3_1_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_0_zpos.txt",net0.n_3_1_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_0_zneg.txt",net0.n_3_1_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_0_xpos.txt",net0.n_3_1_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_0_xneg.txt",net0.n_3_1_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_0_ypos.txt",net0.n_3_1_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_0_yneg.txt",net0.n_3_1_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_0_zpos.txt",net0.n_3_1_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_0_zneg.txt",net0.n_3_1_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_1_local.txt",net0.n_3_1_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_1_xpos.txt",net0.n_3_1_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_1_xneg.txt",net0.n_3_1_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_1_ypos.txt",net0.n_3_1_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_1_yneg.txt",net0.n_3_1_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_1_zpos.txt",net0.n_3_1_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_1_zneg.txt",net0.n_3_1_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_1_xpos.txt",net0.n_3_1_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_1_xneg.txt",net0.n_3_1_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_1_ypos.txt",net0.n_3_1_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_1_yneg.txt",net0.n_3_1_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_1_zpos.txt",net0.n_3_1_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_1_zneg.txt",net0.n_3_1_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_1_xpos.txt",net0.n_3_1_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_1_xneg.txt",net0.n_3_1_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_1_ypos.txt",net0.n_3_1_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_1_yneg.txt",net0.n_3_1_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_1_zpos.txt",net0.n_3_1_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_1_zneg.txt",net0.n_3_1_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_2_local.txt",net0.n_3_1_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_2_xpos.txt",net0.n_3_1_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_2_xneg.txt",net0.n_3_1_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_2_ypos.txt",net0.n_3_1_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_2_yneg.txt",net0.n_3_1_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_2_zpos.txt",net0.n_3_1_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_2_zneg.txt",net0.n_3_1_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_2_xpos.txt",net0.n_3_1_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_2_xneg.txt",net0.n_3_1_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_2_ypos.txt",net0.n_3_1_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_2_yneg.txt",net0.n_3_1_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_2_zpos.txt",net0.n_3_1_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_2_zneg.txt",net0.n_3_1_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_2_xpos.txt",net0.n_3_1_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_2_xneg.txt",net0.n_3_1_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_2_ypos.txt",net0.n_3_1_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_2_yneg.txt",net0.n_3_1_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_2_zpos.txt",net0.n_3_1_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_2_zneg.txt",net0.n_3_1_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_3_local.txt",net0.n_3_1_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_3_xpos.txt",net0.n_3_1_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_3_xneg.txt",net0.n_3_1_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_3_ypos.txt",net0.n_3_1_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_3_yneg.txt",net0.n_3_1_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_3_zpos.txt",net0.n_3_1_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_3_zneg.txt",net0.n_3_1_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_3_xpos.txt",net0.n_3_1_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_3_xneg.txt",net0.n_3_1_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_3_ypos.txt",net0.n_3_1_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_3_yneg.txt",net0.n_3_1_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_3_zpos.txt",net0.n_3_1_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_3_zneg.txt",net0.n_3_1_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_3_xpos.txt",net0.n_3_1_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_3_xneg.txt",net0.n_3_1_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_3_ypos.txt",net0.n_3_1_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_3_yneg.txt",net0.n_3_1_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_3_zpos.txt",net0.n_3_1_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_3_zneg.txt",net0.n_3_1_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_4_local.txt",net0.n_3_1_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_4_xpos.txt",net0.n_3_1_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_4_xneg.txt",net0.n_3_1_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_4_ypos.txt",net0.n_3_1_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_4_yneg.txt",net0.n_3_1_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_4_zpos.txt",net0.n_3_1_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_4_zneg.txt",net0.n_3_1_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_4_xpos.txt",net0.n_3_1_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_4_xneg.txt",net0.n_3_1_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_4_ypos.txt",net0.n_3_1_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_4_yneg.txt",net0.n_3_1_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_4_zpos.txt",net0.n_3_1_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_4_zneg.txt",net0.n_3_1_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_4_xpos.txt",net0.n_3_1_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_4_xneg.txt",net0.n_3_1_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_4_ypos.txt",net0.n_3_1_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_4_yneg.txt",net0.n_3_1_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_4_zpos.txt",net0.n_3_1_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_4_zneg.txt",net0.n_3_1_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_5_local.txt",net0.n_3_1_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_5_xpos.txt",net0.n_3_1_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_5_xneg.txt",net0.n_3_1_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_5_ypos.txt",net0.n_3_1_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_5_yneg.txt",net0.n_3_1_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_5_zpos.txt",net0.n_3_1_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_5_zneg.txt",net0.n_3_1_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_5_xpos.txt",net0.n_3_1_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_5_xneg.txt",net0.n_3_1_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_5_ypos.txt",net0.n_3_1_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_5_yneg.txt",net0.n_3_1_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_5_zpos.txt",net0.n_3_1_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_5_zneg.txt",net0.n_3_1_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_5_xpos.txt",net0.n_3_1_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_5_xneg.txt",net0.n_3_1_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_5_ypos.txt",net0.n_3_1_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_5_yneg.txt",net0.n_3_1_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_5_zpos.txt",net0.n_3_1_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_5_zneg.txt",net0.n_3_1_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_6_local.txt",net0.n_3_1_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_6_xpos.txt",net0.n_3_1_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_6_xneg.txt",net0.n_3_1_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_6_ypos.txt",net0.n_3_1_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_6_yneg.txt",net0.n_3_1_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_6_zpos.txt",net0.n_3_1_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_6_zneg.txt",net0.n_3_1_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_6_xpos.txt",net0.n_3_1_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_6_xneg.txt",net0.n_3_1_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_6_ypos.txt",net0.n_3_1_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_6_yneg.txt",net0.n_3_1_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_6_zpos.txt",net0.n_3_1_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_6_zneg.txt",net0.n_3_1_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_6_xpos.txt",net0.n_3_1_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_6_xneg.txt",net0.n_3_1_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_6_ypos.txt",net0.n_3_1_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_6_yneg.txt",net0.n_3_1_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_6_zpos.txt",net0.n_3_1_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_6_zneg.txt",net0.n_3_1_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_7_local.txt",net0.n_3_1_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_7_xpos.txt",net0.n_3_1_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_7_xneg.txt",net0.n_3_1_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_7_ypos.txt",net0.n_3_1_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_7_yneg.txt",net0.n_3_1_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_7_zpos.txt",net0.n_3_1_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_1_7_zneg.txt",net0.n_3_1_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_7_xpos.txt",net0.n_3_1_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_7_xneg.txt",net0.n_3_1_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_7_ypos.txt",net0.n_3_1_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_7_yneg.txt",net0.n_3_1_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_7_zpos.txt",net0.n_3_1_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_1_7_zneg.txt",net0.n_3_1_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_7_xpos.txt",net0.n_3_1_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_7_xneg.txt",net0.n_3_1_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_7_ypos.txt",net0.n_3_1_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_7_yneg.txt",net0.n_3_1_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_7_zpos.txt",net0.n_3_1_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_1_7_zneg.txt",net0.n_3_1_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_0_local.txt",net0.n_3_2_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_0_xpos.txt",net0.n_3_2_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_0_xneg.txt",net0.n_3_2_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_0_ypos.txt",net0.n_3_2_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_0_yneg.txt",net0.n_3_2_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_0_zpos.txt",net0.n_3_2_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_0_zneg.txt",net0.n_3_2_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_0_xpos.txt",net0.n_3_2_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_0_xneg.txt",net0.n_3_2_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_0_ypos.txt",net0.n_3_2_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_0_yneg.txt",net0.n_3_2_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_0_zpos.txt",net0.n_3_2_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_0_zneg.txt",net0.n_3_2_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_0_xpos.txt",net0.n_3_2_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_0_xneg.txt",net0.n_3_2_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_0_ypos.txt",net0.n_3_2_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_0_yneg.txt",net0.n_3_2_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_0_zpos.txt",net0.n_3_2_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_0_zneg.txt",net0.n_3_2_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_1_local.txt",net0.n_3_2_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_1_xpos.txt",net0.n_3_2_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_1_xneg.txt",net0.n_3_2_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_1_ypos.txt",net0.n_3_2_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_1_yneg.txt",net0.n_3_2_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_1_zpos.txt",net0.n_3_2_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_1_zneg.txt",net0.n_3_2_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_1_xpos.txt",net0.n_3_2_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_1_xneg.txt",net0.n_3_2_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_1_ypos.txt",net0.n_3_2_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_1_yneg.txt",net0.n_3_2_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_1_zpos.txt",net0.n_3_2_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_1_zneg.txt",net0.n_3_2_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_1_xpos.txt",net0.n_3_2_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_1_xneg.txt",net0.n_3_2_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_1_ypos.txt",net0.n_3_2_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_1_yneg.txt",net0.n_3_2_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_1_zpos.txt",net0.n_3_2_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_1_zneg.txt",net0.n_3_2_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_2_local.txt",net0.n_3_2_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_2_xpos.txt",net0.n_3_2_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_2_xneg.txt",net0.n_3_2_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_2_ypos.txt",net0.n_3_2_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_2_yneg.txt",net0.n_3_2_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_2_zpos.txt",net0.n_3_2_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_2_zneg.txt",net0.n_3_2_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_2_xpos.txt",net0.n_3_2_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_2_xneg.txt",net0.n_3_2_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_2_ypos.txt",net0.n_3_2_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_2_yneg.txt",net0.n_3_2_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_2_zpos.txt",net0.n_3_2_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_2_zneg.txt",net0.n_3_2_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_2_xpos.txt",net0.n_3_2_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_2_xneg.txt",net0.n_3_2_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_2_ypos.txt",net0.n_3_2_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_2_yneg.txt",net0.n_3_2_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_2_zpos.txt",net0.n_3_2_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_2_zneg.txt",net0.n_3_2_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_3_local.txt",net0.n_3_2_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_3_xpos.txt",net0.n_3_2_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_3_xneg.txt",net0.n_3_2_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_3_ypos.txt",net0.n_3_2_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_3_yneg.txt",net0.n_3_2_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_3_zpos.txt",net0.n_3_2_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_3_zneg.txt",net0.n_3_2_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_3_xpos.txt",net0.n_3_2_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_3_xneg.txt",net0.n_3_2_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_3_ypos.txt",net0.n_3_2_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_3_yneg.txt",net0.n_3_2_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_3_zpos.txt",net0.n_3_2_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_3_zneg.txt",net0.n_3_2_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_3_xpos.txt",net0.n_3_2_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_3_xneg.txt",net0.n_3_2_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_3_ypos.txt",net0.n_3_2_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_3_yneg.txt",net0.n_3_2_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_3_zpos.txt",net0.n_3_2_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_3_zneg.txt",net0.n_3_2_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_4_local.txt",net0.n_3_2_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_4_xpos.txt",net0.n_3_2_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_4_xneg.txt",net0.n_3_2_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_4_ypos.txt",net0.n_3_2_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_4_yneg.txt",net0.n_3_2_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_4_zpos.txt",net0.n_3_2_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_4_zneg.txt",net0.n_3_2_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_4_xpos.txt",net0.n_3_2_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_4_xneg.txt",net0.n_3_2_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_4_ypos.txt",net0.n_3_2_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_4_yneg.txt",net0.n_3_2_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_4_zpos.txt",net0.n_3_2_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_4_zneg.txt",net0.n_3_2_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_4_xpos.txt",net0.n_3_2_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_4_xneg.txt",net0.n_3_2_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_4_ypos.txt",net0.n_3_2_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_4_yneg.txt",net0.n_3_2_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_4_zpos.txt",net0.n_3_2_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_4_zneg.txt",net0.n_3_2_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_5_local.txt",net0.n_3_2_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_5_xpos.txt",net0.n_3_2_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_5_xneg.txt",net0.n_3_2_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_5_ypos.txt",net0.n_3_2_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_5_yneg.txt",net0.n_3_2_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_5_zpos.txt",net0.n_3_2_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_5_zneg.txt",net0.n_3_2_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_5_xpos.txt",net0.n_3_2_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_5_xneg.txt",net0.n_3_2_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_5_ypos.txt",net0.n_3_2_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_5_yneg.txt",net0.n_3_2_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_5_zpos.txt",net0.n_3_2_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_5_zneg.txt",net0.n_3_2_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_5_xpos.txt",net0.n_3_2_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_5_xneg.txt",net0.n_3_2_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_5_ypos.txt",net0.n_3_2_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_5_yneg.txt",net0.n_3_2_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_5_zpos.txt",net0.n_3_2_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_5_zneg.txt",net0.n_3_2_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_6_local.txt",net0.n_3_2_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_6_xpos.txt",net0.n_3_2_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_6_xneg.txt",net0.n_3_2_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_6_ypos.txt",net0.n_3_2_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_6_yneg.txt",net0.n_3_2_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_6_zpos.txt",net0.n_3_2_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_6_zneg.txt",net0.n_3_2_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_6_xpos.txt",net0.n_3_2_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_6_xneg.txt",net0.n_3_2_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_6_ypos.txt",net0.n_3_2_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_6_yneg.txt",net0.n_3_2_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_6_zpos.txt",net0.n_3_2_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_6_zneg.txt",net0.n_3_2_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_6_xpos.txt",net0.n_3_2_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_6_xneg.txt",net0.n_3_2_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_6_ypos.txt",net0.n_3_2_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_6_yneg.txt",net0.n_3_2_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_6_zpos.txt",net0.n_3_2_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_6_zneg.txt",net0.n_3_2_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_7_local.txt",net0.n_3_2_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_7_xpos.txt",net0.n_3_2_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_7_xneg.txt",net0.n_3_2_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_7_ypos.txt",net0.n_3_2_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_7_yneg.txt",net0.n_3_2_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_7_zpos.txt",net0.n_3_2_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_2_7_zneg.txt",net0.n_3_2_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_7_xpos.txt",net0.n_3_2_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_7_xneg.txt",net0.n_3_2_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_7_ypos.txt",net0.n_3_2_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_7_yneg.txt",net0.n_3_2_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_7_zpos.txt",net0.n_3_2_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_2_7_zneg.txt",net0.n_3_2_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_7_xpos.txt",net0.n_3_2_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_7_xneg.txt",net0.n_3_2_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_7_ypos.txt",net0.n_3_2_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_7_yneg.txt",net0.n_3_2_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_7_zpos.txt",net0.n_3_2_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_2_7_zneg.txt",net0.n_3_2_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_0_local.txt",net0.n_3_3_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_0_xpos.txt",net0.n_3_3_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_0_xneg.txt",net0.n_3_3_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_0_ypos.txt",net0.n_3_3_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_0_yneg.txt",net0.n_3_3_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_0_zpos.txt",net0.n_3_3_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_0_zneg.txt",net0.n_3_3_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_0_xpos.txt",net0.n_3_3_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_0_xneg.txt",net0.n_3_3_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_0_ypos.txt",net0.n_3_3_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_0_yneg.txt",net0.n_3_3_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_0_zpos.txt",net0.n_3_3_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_0_zneg.txt",net0.n_3_3_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_0_xpos.txt",net0.n_3_3_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_0_xneg.txt",net0.n_3_3_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_0_ypos.txt",net0.n_3_3_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_0_yneg.txt",net0.n_3_3_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_0_zpos.txt",net0.n_3_3_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_0_zneg.txt",net0.n_3_3_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_1_local.txt",net0.n_3_3_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_1_xpos.txt",net0.n_3_3_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_1_xneg.txt",net0.n_3_3_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_1_ypos.txt",net0.n_3_3_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_1_yneg.txt",net0.n_3_3_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_1_zpos.txt",net0.n_3_3_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_1_zneg.txt",net0.n_3_3_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_1_xpos.txt",net0.n_3_3_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_1_xneg.txt",net0.n_3_3_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_1_ypos.txt",net0.n_3_3_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_1_yneg.txt",net0.n_3_3_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_1_zpos.txt",net0.n_3_3_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_1_zneg.txt",net0.n_3_3_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_1_xpos.txt",net0.n_3_3_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_1_xneg.txt",net0.n_3_3_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_1_ypos.txt",net0.n_3_3_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_1_yneg.txt",net0.n_3_3_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_1_zpos.txt",net0.n_3_3_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_1_zneg.txt",net0.n_3_3_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_2_local.txt",net0.n_3_3_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_2_xpos.txt",net0.n_3_3_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_2_xneg.txt",net0.n_3_3_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_2_ypos.txt",net0.n_3_3_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_2_yneg.txt",net0.n_3_3_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_2_zpos.txt",net0.n_3_3_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_2_zneg.txt",net0.n_3_3_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_2_xpos.txt",net0.n_3_3_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_2_xneg.txt",net0.n_3_3_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_2_ypos.txt",net0.n_3_3_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_2_yneg.txt",net0.n_3_3_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_2_zpos.txt",net0.n_3_3_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_2_zneg.txt",net0.n_3_3_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_2_xpos.txt",net0.n_3_3_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_2_xneg.txt",net0.n_3_3_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_2_ypos.txt",net0.n_3_3_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_2_yneg.txt",net0.n_3_3_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_2_zpos.txt",net0.n_3_3_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_2_zneg.txt",net0.n_3_3_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_3_local.txt",net0.n_3_3_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_3_xpos.txt",net0.n_3_3_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_3_xneg.txt",net0.n_3_3_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_3_ypos.txt",net0.n_3_3_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_3_yneg.txt",net0.n_3_3_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_3_zpos.txt",net0.n_3_3_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_3_zneg.txt",net0.n_3_3_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_3_xpos.txt",net0.n_3_3_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_3_xneg.txt",net0.n_3_3_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_3_ypos.txt",net0.n_3_3_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_3_yneg.txt",net0.n_3_3_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_3_zpos.txt",net0.n_3_3_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_3_zneg.txt",net0.n_3_3_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_3_xpos.txt",net0.n_3_3_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_3_xneg.txt",net0.n_3_3_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_3_ypos.txt",net0.n_3_3_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_3_yneg.txt",net0.n_3_3_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_3_zpos.txt",net0.n_3_3_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_3_zneg.txt",net0.n_3_3_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_4_local.txt",net0.n_3_3_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_4_xpos.txt",net0.n_3_3_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_4_xneg.txt",net0.n_3_3_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_4_ypos.txt",net0.n_3_3_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_4_yneg.txt",net0.n_3_3_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_4_zpos.txt",net0.n_3_3_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_4_zneg.txt",net0.n_3_3_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_4_xpos.txt",net0.n_3_3_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_4_xneg.txt",net0.n_3_3_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_4_ypos.txt",net0.n_3_3_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_4_yneg.txt",net0.n_3_3_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_4_zpos.txt",net0.n_3_3_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_4_zneg.txt",net0.n_3_3_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_4_xpos.txt",net0.n_3_3_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_4_xneg.txt",net0.n_3_3_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_4_ypos.txt",net0.n_3_3_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_4_yneg.txt",net0.n_3_3_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_4_zpos.txt",net0.n_3_3_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_4_zneg.txt",net0.n_3_3_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_5_local.txt",net0.n_3_3_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_5_xpos.txt",net0.n_3_3_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_5_xneg.txt",net0.n_3_3_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_5_ypos.txt",net0.n_3_3_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_5_yneg.txt",net0.n_3_3_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_5_zpos.txt",net0.n_3_3_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_5_zneg.txt",net0.n_3_3_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_5_xpos.txt",net0.n_3_3_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_5_xneg.txt",net0.n_3_3_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_5_ypos.txt",net0.n_3_3_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_5_yneg.txt",net0.n_3_3_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_5_zpos.txt",net0.n_3_3_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_5_zneg.txt",net0.n_3_3_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_5_xpos.txt",net0.n_3_3_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_5_xneg.txt",net0.n_3_3_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_5_ypos.txt",net0.n_3_3_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_5_yneg.txt",net0.n_3_3_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_5_zpos.txt",net0.n_3_3_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_5_zneg.txt",net0.n_3_3_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_6_local.txt",net0.n_3_3_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_6_xpos.txt",net0.n_3_3_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_6_xneg.txt",net0.n_3_3_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_6_ypos.txt",net0.n_3_3_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_6_yneg.txt",net0.n_3_3_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_6_zpos.txt",net0.n_3_3_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_6_zneg.txt",net0.n_3_3_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_6_xpos.txt",net0.n_3_3_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_6_xneg.txt",net0.n_3_3_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_6_ypos.txt",net0.n_3_3_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_6_yneg.txt",net0.n_3_3_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_6_zpos.txt",net0.n_3_3_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_6_zneg.txt",net0.n_3_3_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_6_xpos.txt",net0.n_3_3_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_6_xneg.txt",net0.n_3_3_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_6_ypos.txt",net0.n_3_3_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_6_yneg.txt",net0.n_3_3_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_6_zpos.txt",net0.n_3_3_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_6_zneg.txt",net0.n_3_3_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_7_local.txt",net0.n_3_3_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_7_xpos.txt",net0.n_3_3_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_7_xneg.txt",net0.n_3_3_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_7_ypos.txt",net0.n_3_3_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_7_yneg.txt",net0.n_3_3_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_7_zpos.txt",net0.n_3_3_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_3_7_zneg.txt",net0.n_3_3_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_7_xpos.txt",net0.n_3_3_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_7_xneg.txt",net0.n_3_3_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_7_ypos.txt",net0.n_3_3_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_7_yneg.txt",net0.n_3_3_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_7_zpos.txt",net0.n_3_3_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_3_7_zneg.txt",net0.n_3_3_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_7_xpos.txt",net0.n_3_3_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_7_xneg.txt",net0.n_3_3_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_7_ypos.txt",net0.n_3_3_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_7_yneg.txt",net0.n_3_3_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_7_zpos.txt",net0.n_3_3_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_3_7_zneg.txt",net0.n_3_3_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_0_local.txt",net0.n_3_4_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_0_xpos.txt",net0.n_3_4_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_0_xneg.txt",net0.n_3_4_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_0_ypos.txt",net0.n_3_4_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_0_yneg.txt",net0.n_3_4_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_0_zpos.txt",net0.n_3_4_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_0_zneg.txt",net0.n_3_4_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_0_xpos.txt",net0.n_3_4_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_0_xneg.txt",net0.n_3_4_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_0_ypos.txt",net0.n_3_4_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_0_yneg.txt",net0.n_3_4_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_0_zpos.txt",net0.n_3_4_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_0_zneg.txt",net0.n_3_4_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_0_xpos.txt",net0.n_3_4_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_0_xneg.txt",net0.n_3_4_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_0_ypos.txt",net0.n_3_4_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_0_yneg.txt",net0.n_3_4_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_0_zpos.txt",net0.n_3_4_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_0_zneg.txt",net0.n_3_4_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_1_local.txt",net0.n_3_4_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_1_xpos.txt",net0.n_3_4_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_1_xneg.txt",net0.n_3_4_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_1_ypos.txt",net0.n_3_4_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_1_yneg.txt",net0.n_3_4_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_1_zpos.txt",net0.n_3_4_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_1_zneg.txt",net0.n_3_4_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_1_xpos.txt",net0.n_3_4_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_1_xneg.txt",net0.n_3_4_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_1_ypos.txt",net0.n_3_4_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_1_yneg.txt",net0.n_3_4_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_1_zpos.txt",net0.n_3_4_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_1_zneg.txt",net0.n_3_4_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_1_xpos.txt",net0.n_3_4_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_1_xneg.txt",net0.n_3_4_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_1_ypos.txt",net0.n_3_4_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_1_yneg.txt",net0.n_3_4_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_1_zpos.txt",net0.n_3_4_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_1_zneg.txt",net0.n_3_4_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_2_local.txt",net0.n_3_4_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_2_xpos.txt",net0.n_3_4_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_2_xneg.txt",net0.n_3_4_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_2_ypos.txt",net0.n_3_4_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_2_yneg.txt",net0.n_3_4_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_2_zpos.txt",net0.n_3_4_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_2_zneg.txt",net0.n_3_4_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_2_xpos.txt",net0.n_3_4_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_2_xneg.txt",net0.n_3_4_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_2_ypos.txt",net0.n_3_4_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_2_yneg.txt",net0.n_3_4_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_2_zpos.txt",net0.n_3_4_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_2_zneg.txt",net0.n_3_4_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_2_xpos.txt",net0.n_3_4_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_2_xneg.txt",net0.n_3_4_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_2_ypos.txt",net0.n_3_4_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_2_yneg.txt",net0.n_3_4_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_2_zpos.txt",net0.n_3_4_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_2_zneg.txt",net0.n_3_4_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_3_local.txt",net0.n_3_4_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_3_xpos.txt",net0.n_3_4_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_3_xneg.txt",net0.n_3_4_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_3_ypos.txt",net0.n_3_4_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_3_yneg.txt",net0.n_3_4_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_3_zpos.txt",net0.n_3_4_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_3_zneg.txt",net0.n_3_4_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_3_xpos.txt",net0.n_3_4_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_3_xneg.txt",net0.n_3_4_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_3_ypos.txt",net0.n_3_4_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_3_yneg.txt",net0.n_3_4_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_3_zpos.txt",net0.n_3_4_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_3_zneg.txt",net0.n_3_4_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_3_xpos.txt",net0.n_3_4_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_3_xneg.txt",net0.n_3_4_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_3_ypos.txt",net0.n_3_4_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_3_yneg.txt",net0.n_3_4_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_3_zpos.txt",net0.n_3_4_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_3_zneg.txt",net0.n_3_4_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_4_local.txt",net0.n_3_4_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_4_xpos.txt",net0.n_3_4_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_4_xneg.txt",net0.n_3_4_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_4_ypos.txt",net0.n_3_4_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_4_yneg.txt",net0.n_3_4_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_4_zpos.txt",net0.n_3_4_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_4_zneg.txt",net0.n_3_4_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_4_xpos.txt",net0.n_3_4_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_4_xneg.txt",net0.n_3_4_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_4_ypos.txt",net0.n_3_4_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_4_yneg.txt",net0.n_3_4_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_4_zpos.txt",net0.n_3_4_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_4_zneg.txt",net0.n_3_4_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_4_xpos.txt",net0.n_3_4_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_4_xneg.txt",net0.n_3_4_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_4_ypos.txt",net0.n_3_4_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_4_yneg.txt",net0.n_3_4_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_4_zpos.txt",net0.n_3_4_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_4_zneg.txt",net0.n_3_4_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_5_local.txt",net0.n_3_4_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_5_xpos.txt",net0.n_3_4_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_5_xneg.txt",net0.n_3_4_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_5_ypos.txt",net0.n_3_4_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_5_yneg.txt",net0.n_3_4_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_5_zpos.txt",net0.n_3_4_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_5_zneg.txt",net0.n_3_4_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_5_xpos.txt",net0.n_3_4_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_5_xneg.txt",net0.n_3_4_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_5_ypos.txt",net0.n_3_4_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_5_yneg.txt",net0.n_3_4_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_5_zpos.txt",net0.n_3_4_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_5_zneg.txt",net0.n_3_4_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_5_xpos.txt",net0.n_3_4_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_5_xneg.txt",net0.n_3_4_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_5_ypos.txt",net0.n_3_4_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_5_yneg.txt",net0.n_3_4_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_5_zpos.txt",net0.n_3_4_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_5_zneg.txt",net0.n_3_4_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_6_local.txt",net0.n_3_4_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_6_xpos.txt",net0.n_3_4_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_6_xneg.txt",net0.n_3_4_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_6_ypos.txt",net0.n_3_4_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_6_yneg.txt",net0.n_3_4_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_6_zpos.txt",net0.n_3_4_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_6_zneg.txt",net0.n_3_4_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_6_xpos.txt",net0.n_3_4_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_6_xneg.txt",net0.n_3_4_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_6_ypos.txt",net0.n_3_4_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_6_yneg.txt",net0.n_3_4_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_6_zpos.txt",net0.n_3_4_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_6_zneg.txt",net0.n_3_4_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_6_xpos.txt",net0.n_3_4_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_6_xneg.txt",net0.n_3_4_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_6_ypos.txt",net0.n_3_4_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_6_yneg.txt",net0.n_3_4_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_6_zpos.txt",net0.n_3_4_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_6_zneg.txt",net0.n_3_4_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_7_local.txt",net0.n_3_4_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_7_xpos.txt",net0.n_3_4_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_7_xneg.txt",net0.n_3_4_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_7_ypos.txt",net0.n_3_4_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_7_yneg.txt",net0.n_3_4_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_7_zpos.txt",net0.n_3_4_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_4_7_zneg.txt",net0.n_3_4_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_7_xpos.txt",net0.n_3_4_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_7_xneg.txt",net0.n_3_4_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_7_ypos.txt",net0.n_3_4_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_7_yneg.txt",net0.n_3_4_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_7_zpos.txt",net0.n_3_4_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_4_7_zneg.txt",net0.n_3_4_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_7_xpos.txt",net0.n_3_4_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_7_xneg.txt",net0.n_3_4_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_7_ypos.txt",net0.n_3_4_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_7_yneg.txt",net0.n_3_4_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_7_zpos.txt",net0.n_3_4_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_4_7_zneg.txt",net0.n_3_4_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_0_local.txt",net0.n_3_5_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_0_xpos.txt",net0.n_3_5_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_0_xneg.txt",net0.n_3_5_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_0_ypos.txt",net0.n_3_5_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_0_yneg.txt",net0.n_3_5_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_0_zpos.txt",net0.n_3_5_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_0_zneg.txt",net0.n_3_5_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_0_xpos.txt",net0.n_3_5_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_0_xneg.txt",net0.n_3_5_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_0_ypos.txt",net0.n_3_5_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_0_yneg.txt",net0.n_3_5_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_0_zpos.txt",net0.n_3_5_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_0_zneg.txt",net0.n_3_5_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_0_xpos.txt",net0.n_3_5_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_0_xneg.txt",net0.n_3_5_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_0_ypos.txt",net0.n_3_5_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_0_yneg.txt",net0.n_3_5_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_0_zpos.txt",net0.n_3_5_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_0_zneg.txt",net0.n_3_5_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_1_local.txt",net0.n_3_5_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_1_xpos.txt",net0.n_3_5_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_1_xneg.txt",net0.n_3_5_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_1_ypos.txt",net0.n_3_5_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_1_yneg.txt",net0.n_3_5_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_1_zpos.txt",net0.n_3_5_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_1_zneg.txt",net0.n_3_5_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_1_xpos.txt",net0.n_3_5_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_1_xneg.txt",net0.n_3_5_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_1_ypos.txt",net0.n_3_5_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_1_yneg.txt",net0.n_3_5_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_1_zpos.txt",net0.n_3_5_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_1_zneg.txt",net0.n_3_5_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_1_xpos.txt",net0.n_3_5_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_1_xneg.txt",net0.n_3_5_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_1_ypos.txt",net0.n_3_5_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_1_yneg.txt",net0.n_3_5_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_1_zpos.txt",net0.n_3_5_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_1_zneg.txt",net0.n_3_5_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_2_local.txt",net0.n_3_5_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_2_xpos.txt",net0.n_3_5_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_2_xneg.txt",net0.n_3_5_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_2_ypos.txt",net0.n_3_5_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_2_yneg.txt",net0.n_3_5_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_2_zpos.txt",net0.n_3_5_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_2_zneg.txt",net0.n_3_5_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_2_xpos.txt",net0.n_3_5_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_2_xneg.txt",net0.n_3_5_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_2_ypos.txt",net0.n_3_5_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_2_yneg.txt",net0.n_3_5_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_2_zpos.txt",net0.n_3_5_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_2_zneg.txt",net0.n_3_5_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_2_xpos.txt",net0.n_3_5_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_2_xneg.txt",net0.n_3_5_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_2_ypos.txt",net0.n_3_5_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_2_yneg.txt",net0.n_3_5_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_2_zpos.txt",net0.n_3_5_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_2_zneg.txt",net0.n_3_5_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_3_local.txt",net0.n_3_5_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_3_xpos.txt",net0.n_3_5_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_3_xneg.txt",net0.n_3_5_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_3_ypos.txt",net0.n_3_5_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_3_yneg.txt",net0.n_3_5_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_3_zpos.txt",net0.n_3_5_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_3_zneg.txt",net0.n_3_5_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_3_xpos.txt",net0.n_3_5_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_3_xneg.txt",net0.n_3_5_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_3_ypos.txt",net0.n_3_5_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_3_yneg.txt",net0.n_3_5_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_3_zpos.txt",net0.n_3_5_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_3_zneg.txt",net0.n_3_5_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_3_xpos.txt",net0.n_3_5_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_3_xneg.txt",net0.n_3_5_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_3_ypos.txt",net0.n_3_5_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_3_yneg.txt",net0.n_3_5_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_3_zpos.txt",net0.n_3_5_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_3_zneg.txt",net0.n_3_5_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_4_local.txt",net0.n_3_5_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_4_xpos.txt",net0.n_3_5_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_4_xneg.txt",net0.n_3_5_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_4_ypos.txt",net0.n_3_5_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_4_yneg.txt",net0.n_3_5_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_4_zpos.txt",net0.n_3_5_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_4_zneg.txt",net0.n_3_5_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_4_xpos.txt",net0.n_3_5_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_4_xneg.txt",net0.n_3_5_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_4_ypos.txt",net0.n_3_5_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_4_yneg.txt",net0.n_3_5_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_4_zpos.txt",net0.n_3_5_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_4_zneg.txt",net0.n_3_5_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_4_xpos.txt",net0.n_3_5_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_4_xneg.txt",net0.n_3_5_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_4_ypos.txt",net0.n_3_5_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_4_yneg.txt",net0.n_3_5_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_4_zpos.txt",net0.n_3_5_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_4_zneg.txt",net0.n_3_5_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_5_local.txt",net0.n_3_5_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_5_xpos.txt",net0.n_3_5_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_5_xneg.txt",net0.n_3_5_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_5_ypos.txt",net0.n_3_5_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_5_yneg.txt",net0.n_3_5_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_5_zpos.txt",net0.n_3_5_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_5_zneg.txt",net0.n_3_5_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_5_xpos.txt",net0.n_3_5_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_5_xneg.txt",net0.n_3_5_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_5_ypos.txt",net0.n_3_5_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_5_yneg.txt",net0.n_3_5_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_5_zpos.txt",net0.n_3_5_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_5_zneg.txt",net0.n_3_5_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_5_xpos.txt",net0.n_3_5_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_5_xneg.txt",net0.n_3_5_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_5_ypos.txt",net0.n_3_5_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_5_yneg.txt",net0.n_3_5_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_5_zpos.txt",net0.n_3_5_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_5_zneg.txt",net0.n_3_5_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_6_local.txt",net0.n_3_5_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_6_xpos.txt",net0.n_3_5_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_6_xneg.txt",net0.n_3_5_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_6_ypos.txt",net0.n_3_5_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_6_yneg.txt",net0.n_3_5_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_6_zpos.txt",net0.n_3_5_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_6_zneg.txt",net0.n_3_5_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_6_xpos.txt",net0.n_3_5_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_6_xneg.txt",net0.n_3_5_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_6_ypos.txt",net0.n_3_5_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_6_yneg.txt",net0.n_3_5_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_6_zpos.txt",net0.n_3_5_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_6_zneg.txt",net0.n_3_5_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_6_xpos.txt",net0.n_3_5_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_6_xneg.txt",net0.n_3_5_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_6_ypos.txt",net0.n_3_5_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_6_yneg.txt",net0.n_3_5_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_6_zpos.txt",net0.n_3_5_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_6_zneg.txt",net0.n_3_5_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_7_local.txt",net0.n_3_5_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_7_xpos.txt",net0.n_3_5_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_7_xneg.txt",net0.n_3_5_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_7_ypos.txt",net0.n_3_5_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_7_yneg.txt",net0.n_3_5_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_7_zpos.txt",net0.n_3_5_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_5_7_zneg.txt",net0.n_3_5_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_7_xpos.txt",net0.n_3_5_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_7_xneg.txt",net0.n_3_5_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_7_ypos.txt",net0.n_3_5_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_7_yneg.txt",net0.n_3_5_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_7_zpos.txt",net0.n_3_5_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_5_7_zneg.txt",net0.n_3_5_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_7_xpos.txt",net0.n_3_5_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_7_xneg.txt",net0.n_3_5_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_7_ypos.txt",net0.n_3_5_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_7_yneg.txt",net0.n_3_5_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_7_zpos.txt",net0.n_3_5_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_5_7_zneg.txt",net0.n_3_5_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_0_local.txt",net0.n_3_6_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_0_xpos.txt",net0.n_3_6_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_0_xneg.txt",net0.n_3_6_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_0_ypos.txt",net0.n_3_6_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_0_yneg.txt",net0.n_3_6_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_0_zpos.txt",net0.n_3_6_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_0_zneg.txt",net0.n_3_6_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_0_xpos.txt",net0.n_3_6_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_0_xneg.txt",net0.n_3_6_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_0_ypos.txt",net0.n_3_6_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_0_yneg.txt",net0.n_3_6_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_0_zpos.txt",net0.n_3_6_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_0_zneg.txt",net0.n_3_6_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_0_xpos.txt",net0.n_3_6_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_0_xneg.txt",net0.n_3_6_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_0_ypos.txt",net0.n_3_6_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_0_yneg.txt",net0.n_3_6_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_0_zpos.txt",net0.n_3_6_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_0_zneg.txt",net0.n_3_6_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_1_local.txt",net0.n_3_6_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_1_xpos.txt",net0.n_3_6_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_1_xneg.txt",net0.n_3_6_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_1_ypos.txt",net0.n_3_6_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_1_yneg.txt",net0.n_3_6_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_1_zpos.txt",net0.n_3_6_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_1_zneg.txt",net0.n_3_6_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_1_xpos.txt",net0.n_3_6_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_1_xneg.txt",net0.n_3_6_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_1_ypos.txt",net0.n_3_6_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_1_yneg.txt",net0.n_3_6_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_1_zpos.txt",net0.n_3_6_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_1_zneg.txt",net0.n_3_6_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_1_xpos.txt",net0.n_3_6_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_1_xneg.txt",net0.n_3_6_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_1_ypos.txt",net0.n_3_6_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_1_yneg.txt",net0.n_3_6_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_1_zpos.txt",net0.n_3_6_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_1_zneg.txt",net0.n_3_6_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_2_local.txt",net0.n_3_6_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_2_xpos.txt",net0.n_3_6_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_2_xneg.txt",net0.n_3_6_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_2_ypos.txt",net0.n_3_6_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_2_yneg.txt",net0.n_3_6_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_2_zpos.txt",net0.n_3_6_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_2_zneg.txt",net0.n_3_6_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_2_xpos.txt",net0.n_3_6_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_2_xneg.txt",net0.n_3_6_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_2_ypos.txt",net0.n_3_6_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_2_yneg.txt",net0.n_3_6_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_2_zpos.txt",net0.n_3_6_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_2_zneg.txt",net0.n_3_6_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_2_xpos.txt",net0.n_3_6_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_2_xneg.txt",net0.n_3_6_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_2_ypos.txt",net0.n_3_6_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_2_yneg.txt",net0.n_3_6_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_2_zpos.txt",net0.n_3_6_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_2_zneg.txt",net0.n_3_6_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_3_local.txt",net0.n_3_6_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_3_xpos.txt",net0.n_3_6_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_3_xneg.txt",net0.n_3_6_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_3_ypos.txt",net0.n_3_6_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_3_yneg.txt",net0.n_3_6_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_3_zpos.txt",net0.n_3_6_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_3_zneg.txt",net0.n_3_6_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_3_xpos.txt",net0.n_3_6_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_3_xneg.txt",net0.n_3_6_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_3_ypos.txt",net0.n_3_6_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_3_yneg.txt",net0.n_3_6_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_3_zpos.txt",net0.n_3_6_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_3_zneg.txt",net0.n_3_6_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_3_xpos.txt",net0.n_3_6_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_3_xneg.txt",net0.n_3_6_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_3_ypos.txt",net0.n_3_6_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_3_yneg.txt",net0.n_3_6_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_3_zpos.txt",net0.n_3_6_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_3_zneg.txt",net0.n_3_6_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_4_local.txt",net0.n_3_6_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_4_xpos.txt",net0.n_3_6_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_4_xneg.txt",net0.n_3_6_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_4_ypos.txt",net0.n_3_6_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_4_yneg.txt",net0.n_3_6_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_4_zpos.txt",net0.n_3_6_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_4_zneg.txt",net0.n_3_6_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_4_xpos.txt",net0.n_3_6_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_4_xneg.txt",net0.n_3_6_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_4_ypos.txt",net0.n_3_6_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_4_yneg.txt",net0.n_3_6_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_4_zpos.txt",net0.n_3_6_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_4_zneg.txt",net0.n_3_6_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_4_xpos.txt",net0.n_3_6_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_4_xneg.txt",net0.n_3_6_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_4_ypos.txt",net0.n_3_6_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_4_yneg.txt",net0.n_3_6_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_4_zpos.txt",net0.n_3_6_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_4_zneg.txt",net0.n_3_6_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_5_local.txt",net0.n_3_6_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_5_xpos.txt",net0.n_3_6_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_5_xneg.txt",net0.n_3_6_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_5_ypos.txt",net0.n_3_6_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_5_yneg.txt",net0.n_3_6_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_5_zpos.txt",net0.n_3_6_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_5_zneg.txt",net0.n_3_6_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_5_xpos.txt",net0.n_3_6_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_5_xneg.txt",net0.n_3_6_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_5_ypos.txt",net0.n_3_6_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_5_yneg.txt",net0.n_3_6_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_5_zpos.txt",net0.n_3_6_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_5_zneg.txt",net0.n_3_6_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_5_xpos.txt",net0.n_3_6_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_5_xneg.txt",net0.n_3_6_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_5_ypos.txt",net0.n_3_6_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_5_yneg.txt",net0.n_3_6_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_5_zpos.txt",net0.n_3_6_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_5_zneg.txt",net0.n_3_6_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_6_local.txt",net0.n_3_6_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_6_xpos.txt",net0.n_3_6_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_6_xneg.txt",net0.n_3_6_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_6_ypos.txt",net0.n_3_6_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_6_yneg.txt",net0.n_3_6_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_6_zpos.txt",net0.n_3_6_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_6_zneg.txt",net0.n_3_6_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_6_xpos.txt",net0.n_3_6_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_6_xneg.txt",net0.n_3_6_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_6_ypos.txt",net0.n_3_6_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_6_yneg.txt",net0.n_3_6_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_6_zpos.txt",net0.n_3_6_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_6_zneg.txt",net0.n_3_6_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_6_xpos.txt",net0.n_3_6_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_6_xneg.txt",net0.n_3_6_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_6_ypos.txt",net0.n_3_6_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_6_yneg.txt",net0.n_3_6_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_6_zpos.txt",net0.n_3_6_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_6_zneg.txt",net0.n_3_6_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_7_local.txt",net0.n_3_6_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_7_xpos.txt",net0.n_3_6_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_7_xneg.txt",net0.n_3_6_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_7_ypos.txt",net0.n_3_6_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_7_yneg.txt",net0.n_3_6_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_7_zpos.txt",net0.n_3_6_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_6_7_zneg.txt",net0.n_3_6_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_7_xpos.txt",net0.n_3_6_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_7_xneg.txt",net0.n_3_6_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_7_ypos.txt",net0.n_3_6_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_7_yneg.txt",net0.n_3_6_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_7_zpos.txt",net0.n_3_6_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_6_7_zneg.txt",net0.n_3_6_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_7_xpos.txt",net0.n_3_6_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_7_xneg.txt",net0.n_3_6_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_7_ypos.txt",net0.n_3_6_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_7_yneg.txt",net0.n_3_6_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_7_zpos.txt",net0.n_3_6_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_6_7_zneg.txt",net0.n_3_6_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_0_local.txt",net0.n_3_7_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_0_xpos.txt",net0.n_3_7_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_0_xneg.txt",net0.n_3_7_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_0_ypos.txt",net0.n_3_7_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_0_yneg.txt",net0.n_3_7_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_0_zpos.txt",net0.n_3_7_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_0_zneg.txt",net0.n_3_7_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_0_xpos.txt",net0.n_3_7_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_0_xneg.txt",net0.n_3_7_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_0_ypos.txt",net0.n_3_7_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_0_yneg.txt",net0.n_3_7_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_0_zpos.txt",net0.n_3_7_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_0_zneg.txt",net0.n_3_7_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_0_xpos.txt",net0.n_3_7_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_0_xneg.txt",net0.n_3_7_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_0_ypos.txt",net0.n_3_7_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_0_yneg.txt",net0.n_3_7_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_0_zpos.txt",net0.n_3_7_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_0_zneg.txt",net0.n_3_7_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_1_local.txt",net0.n_3_7_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_1_xpos.txt",net0.n_3_7_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_1_xneg.txt",net0.n_3_7_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_1_ypos.txt",net0.n_3_7_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_1_yneg.txt",net0.n_3_7_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_1_zpos.txt",net0.n_3_7_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_1_zneg.txt",net0.n_3_7_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_1_xpos.txt",net0.n_3_7_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_1_xneg.txt",net0.n_3_7_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_1_ypos.txt",net0.n_3_7_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_1_yneg.txt",net0.n_3_7_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_1_zpos.txt",net0.n_3_7_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_1_zneg.txt",net0.n_3_7_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_1_xpos.txt",net0.n_3_7_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_1_xneg.txt",net0.n_3_7_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_1_ypos.txt",net0.n_3_7_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_1_yneg.txt",net0.n_3_7_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_1_zpos.txt",net0.n_3_7_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_1_zneg.txt",net0.n_3_7_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_2_local.txt",net0.n_3_7_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_2_xpos.txt",net0.n_3_7_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_2_xneg.txt",net0.n_3_7_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_2_ypos.txt",net0.n_3_7_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_2_yneg.txt",net0.n_3_7_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_2_zpos.txt",net0.n_3_7_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_2_zneg.txt",net0.n_3_7_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_2_xpos.txt",net0.n_3_7_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_2_xneg.txt",net0.n_3_7_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_2_ypos.txt",net0.n_3_7_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_2_yneg.txt",net0.n_3_7_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_2_zpos.txt",net0.n_3_7_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_2_zneg.txt",net0.n_3_7_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_2_xpos.txt",net0.n_3_7_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_2_xneg.txt",net0.n_3_7_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_2_ypos.txt",net0.n_3_7_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_2_yneg.txt",net0.n_3_7_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_2_zpos.txt",net0.n_3_7_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_2_zneg.txt",net0.n_3_7_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_3_local.txt",net0.n_3_7_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_3_xpos.txt",net0.n_3_7_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_3_xneg.txt",net0.n_3_7_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_3_ypos.txt",net0.n_3_7_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_3_yneg.txt",net0.n_3_7_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_3_zpos.txt",net0.n_3_7_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_3_zneg.txt",net0.n_3_7_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_3_xpos.txt",net0.n_3_7_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_3_xneg.txt",net0.n_3_7_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_3_ypos.txt",net0.n_3_7_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_3_yneg.txt",net0.n_3_7_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_3_zpos.txt",net0.n_3_7_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_3_zneg.txt",net0.n_3_7_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_3_xpos.txt",net0.n_3_7_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_3_xneg.txt",net0.n_3_7_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_3_ypos.txt",net0.n_3_7_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_3_yneg.txt",net0.n_3_7_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_3_zpos.txt",net0.n_3_7_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_3_zneg.txt",net0.n_3_7_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_4_local.txt",net0.n_3_7_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_4_xpos.txt",net0.n_3_7_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_4_xneg.txt",net0.n_3_7_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_4_ypos.txt",net0.n_3_7_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_4_yneg.txt",net0.n_3_7_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_4_zpos.txt",net0.n_3_7_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_4_zneg.txt",net0.n_3_7_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_4_xpos.txt",net0.n_3_7_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_4_xneg.txt",net0.n_3_7_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_4_ypos.txt",net0.n_3_7_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_4_yneg.txt",net0.n_3_7_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_4_zpos.txt",net0.n_3_7_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_4_zneg.txt",net0.n_3_7_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_4_xpos.txt",net0.n_3_7_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_4_xneg.txt",net0.n_3_7_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_4_ypos.txt",net0.n_3_7_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_4_yneg.txt",net0.n_3_7_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_4_zpos.txt",net0.n_3_7_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_4_zneg.txt",net0.n_3_7_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_5_local.txt",net0.n_3_7_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_5_xpos.txt",net0.n_3_7_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_5_xneg.txt",net0.n_3_7_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_5_ypos.txt",net0.n_3_7_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_5_yneg.txt",net0.n_3_7_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_5_zpos.txt",net0.n_3_7_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_5_zneg.txt",net0.n_3_7_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_5_xpos.txt",net0.n_3_7_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_5_xneg.txt",net0.n_3_7_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_5_ypos.txt",net0.n_3_7_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_5_yneg.txt",net0.n_3_7_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_5_zpos.txt",net0.n_3_7_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_5_zneg.txt",net0.n_3_7_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_5_xpos.txt",net0.n_3_7_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_5_xneg.txt",net0.n_3_7_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_5_ypos.txt",net0.n_3_7_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_5_yneg.txt",net0.n_3_7_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_5_zpos.txt",net0.n_3_7_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_5_zneg.txt",net0.n_3_7_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_6_local.txt",net0.n_3_7_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_6_xpos.txt",net0.n_3_7_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_6_xneg.txt",net0.n_3_7_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_6_ypos.txt",net0.n_3_7_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_6_yneg.txt",net0.n_3_7_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_6_zpos.txt",net0.n_3_7_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_6_zneg.txt",net0.n_3_7_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_6_xpos.txt",net0.n_3_7_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_6_xneg.txt",net0.n_3_7_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_6_ypos.txt",net0.n_3_7_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_6_yneg.txt",net0.n_3_7_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_6_zpos.txt",net0.n_3_7_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_6_zneg.txt",net0.n_3_7_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_6_xpos.txt",net0.n_3_7_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_6_xneg.txt",net0.n_3_7_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_6_ypos.txt",net0.n_3_7_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_6_yneg.txt",net0.n_3_7_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_6_zpos.txt",net0.n_3_7_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_6_zneg.txt",net0.n_3_7_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_7_local.txt",net0.n_3_7_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_7_xpos.txt",net0.n_3_7_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_7_xneg.txt",net0.n_3_7_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_7_ypos.txt",net0.n_3_7_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_7_yneg.txt",net0.n_3_7_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_7_zpos.txt",net0.n_3_7_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_3_7_7_zneg.txt",net0.n_3_7_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_7_xpos.txt",net0.n_3_7_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_7_xneg.txt",net0.n_3_7_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_7_ypos.txt",net0.n_3_7_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_7_yneg.txt",net0.n_3_7_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_7_zpos.txt",net0.n_3_7_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_3_7_7_zneg.txt",net0.n_3_7_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_7_xpos.txt",net0.n_3_7_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_7_xneg.txt",net0.n_3_7_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_7_ypos.txt",net0.n_3_7_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_7_yneg.txt",net0.n_3_7_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_7_zpos.txt",net0.n_3_7_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_3_7_7_zneg.txt",net0.n_3_7_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_0_local.txt",net0.n_4_0_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_0_xpos.txt",net0.n_4_0_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_0_xneg.txt",net0.n_4_0_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_0_ypos.txt",net0.n_4_0_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_0_yneg.txt",net0.n_4_0_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_0_zpos.txt",net0.n_4_0_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_0_zneg.txt",net0.n_4_0_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_0_xpos.txt",net0.n_4_0_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_0_xneg.txt",net0.n_4_0_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_0_ypos.txt",net0.n_4_0_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_0_yneg.txt",net0.n_4_0_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_0_zpos.txt",net0.n_4_0_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_0_zneg.txt",net0.n_4_0_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_0_xpos.txt",net0.n_4_0_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_0_xneg.txt",net0.n_4_0_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_0_ypos.txt",net0.n_4_0_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_0_yneg.txt",net0.n_4_0_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_0_zpos.txt",net0.n_4_0_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_0_zneg.txt",net0.n_4_0_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_1_local.txt",net0.n_4_0_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_1_xpos.txt",net0.n_4_0_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_1_xneg.txt",net0.n_4_0_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_1_ypos.txt",net0.n_4_0_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_1_yneg.txt",net0.n_4_0_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_1_zpos.txt",net0.n_4_0_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_1_zneg.txt",net0.n_4_0_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_1_xpos.txt",net0.n_4_0_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_1_xneg.txt",net0.n_4_0_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_1_ypos.txt",net0.n_4_0_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_1_yneg.txt",net0.n_4_0_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_1_zpos.txt",net0.n_4_0_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_1_zneg.txt",net0.n_4_0_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_1_xpos.txt",net0.n_4_0_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_1_xneg.txt",net0.n_4_0_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_1_ypos.txt",net0.n_4_0_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_1_yneg.txt",net0.n_4_0_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_1_zpos.txt",net0.n_4_0_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_1_zneg.txt",net0.n_4_0_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_2_local.txt",net0.n_4_0_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_2_xpos.txt",net0.n_4_0_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_2_xneg.txt",net0.n_4_0_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_2_ypos.txt",net0.n_4_0_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_2_yneg.txt",net0.n_4_0_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_2_zpos.txt",net0.n_4_0_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_2_zneg.txt",net0.n_4_0_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_2_xpos.txt",net0.n_4_0_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_2_xneg.txt",net0.n_4_0_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_2_ypos.txt",net0.n_4_0_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_2_yneg.txt",net0.n_4_0_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_2_zpos.txt",net0.n_4_0_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_2_zneg.txt",net0.n_4_0_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_2_xpos.txt",net0.n_4_0_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_2_xneg.txt",net0.n_4_0_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_2_ypos.txt",net0.n_4_0_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_2_yneg.txt",net0.n_4_0_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_2_zpos.txt",net0.n_4_0_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_2_zneg.txt",net0.n_4_0_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_3_local.txt",net0.n_4_0_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_3_xpos.txt",net0.n_4_0_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_3_xneg.txt",net0.n_4_0_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_3_ypos.txt",net0.n_4_0_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_3_yneg.txt",net0.n_4_0_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_3_zpos.txt",net0.n_4_0_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_3_zneg.txt",net0.n_4_0_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_3_xpos.txt",net0.n_4_0_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_3_xneg.txt",net0.n_4_0_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_3_ypos.txt",net0.n_4_0_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_3_yneg.txt",net0.n_4_0_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_3_zpos.txt",net0.n_4_0_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_3_zneg.txt",net0.n_4_0_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_3_xpos.txt",net0.n_4_0_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_3_xneg.txt",net0.n_4_0_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_3_ypos.txt",net0.n_4_0_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_3_yneg.txt",net0.n_4_0_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_3_zpos.txt",net0.n_4_0_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_3_zneg.txt",net0.n_4_0_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_4_local.txt",net0.n_4_0_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_4_xpos.txt",net0.n_4_0_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_4_xneg.txt",net0.n_4_0_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_4_ypos.txt",net0.n_4_0_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_4_yneg.txt",net0.n_4_0_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_4_zpos.txt",net0.n_4_0_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_4_zneg.txt",net0.n_4_0_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_4_xpos.txt",net0.n_4_0_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_4_xneg.txt",net0.n_4_0_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_4_ypos.txt",net0.n_4_0_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_4_yneg.txt",net0.n_4_0_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_4_zpos.txt",net0.n_4_0_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_4_zneg.txt",net0.n_4_0_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_4_xpos.txt",net0.n_4_0_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_4_xneg.txt",net0.n_4_0_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_4_ypos.txt",net0.n_4_0_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_4_yneg.txt",net0.n_4_0_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_4_zpos.txt",net0.n_4_0_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_4_zneg.txt",net0.n_4_0_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_5_local.txt",net0.n_4_0_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_5_xpos.txt",net0.n_4_0_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_5_xneg.txt",net0.n_4_0_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_5_ypos.txt",net0.n_4_0_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_5_yneg.txt",net0.n_4_0_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_5_zpos.txt",net0.n_4_0_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_5_zneg.txt",net0.n_4_0_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_5_xpos.txt",net0.n_4_0_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_5_xneg.txt",net0.n_4_0_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_5_ypos.txt",net0.n_4_0_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_5_yneg.txt",net0.n_4_0_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_5_zpos.txt",net0.n_4_0_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_5_zneg.txt",net0.n_4_0_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_5_xpos.txt",net0.n_4_0_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_5_xneg.txt",net0.n_4_0_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_5_ypos.txt",net0.n_4_0_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_5_yneg.txt",net0.n_4_0_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_5_zpos.txt",net0.n_4_0_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_5_zneg.txt",net0.n_4_0_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_6_local.txt",net0.n_4_0_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_6_xpos.txt",net0.n_4_0_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_6_xneg.txt",net0.n_4_0_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_6_ypos.txt",net0.n_4_0_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_6_yneg.txt",net0.n_4_0_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_6_zpos.txt",net0.n_4_0_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_6_zneg.txt",net0.n_4_0_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_6_xpos.txt",net0.n_4_0_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_6_xneg.txt",net0.n_4_0_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_6_ypos.txt",net0.n_4_0_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_6_yneg.txt",net0.n_4_0_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_6_zpos.txt",net0.n_4_0_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_6_zneg.txt",net0.n_4_0_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_6_xpos.txt",net0.n_4_0_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_6_xneg.txt",net0.n_4_0_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_6_ypos.txt",net0.n_4_0_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_6_yneg.txt",net0.n_4_0_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_6_zpos.txt",net0.n_4_0_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_6_zneg.txt",net0.n_4_0_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_7_local.txt",net0.n_4_0_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_7_xpos.txt",net0.n_4_0_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_7_xneg.txt",net0.n_4_0_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_7_ypos.txt",net0.n_4_0_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_7_yneg.txt",net0.n_4_0_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_7_zpos.txt",net0.n_4_0_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_0_7_zneg.txt",net0.n_4_0_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_7_xpos.txt",net0.n_4_0_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_7_xneg.txt",net0.n_4_0_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_7_ypos.txt",net0.n_4_0_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_7_yneg.txt",net0.n_4_0_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_7_zpos.txt",net0.n_4_0_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_0_7_zneg.txt",net0.n_4_0_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_7_xpos.txt",net0.n_4_0_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_7_xneg.txt",net0.n_4_0_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_7_ypos.txt",net0.n_4_0_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_7_yneg.txt",net0.n_4_0_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_7_zpos.txt",net0.n_4_0_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_0_7_zneg.txt",net0.n_4_0_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_0_local.txt",net0.n_4_1_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_0_xpos.txt",net0.n_4_1_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_0_xneg.txt",net0.n_4_1_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_0_ypos.txt",net0.n_4_1_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_0_yneg.txt",net0.n_4_1_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_0_zpos.txt",net0.n_4_1_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_0_zneg.txt",net0.n_4_1_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_0_xpos.txt",net0.n_4_1_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_0_xneg.txt",net0.n_4_1_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_0_ypos.txt",net0.n_4_1_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_0_yneg.txt",net0.n_4_1_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_0_zpos.txt",net0.n_4_1_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_0_zneg.txt",net0.n_4_1_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_0_xpos.txt",net0.n_4_1_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_0_xneg.txt",net0.n_4_1_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_0_ypos.txt",net0.n_4_1_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_0_yneg.txt",net0.n_4_1_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_0_zpos.txt",net0.n_4_1_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_0_zneg.txt",net0.n_4_1_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_1_local.txt",net0.n_4_1_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_1_xpos.txt",net0.n_4_1_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_1_xneg.txt",net0.n_4_1_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_1_ypos.txt",net0.n_4_1_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_1_yneg.txt",net0.n_4_1_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_1_zpos.txt",net0.n_4_1_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_1_zneg.txt",net0.n_4_1_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_1_xpos.txt",net0.n_4_1_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_1_xneg.txt",net0.n_4_1_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_1_ypos.txt",net0.n_4_1_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_1_yneg.txt",net0.n_4_1_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_1_zpos.txt",net0.n_4_1_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_1_zneg.txt",net0.n_4_1_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_1_xpos.txt",net0.n_4_1_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_1_xneg.txt",net0.n_4_1_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_1_ypos.txt",net0.n_4_1_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_1_yneg.txt",net0.n_4_1_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_1_zpos.txt",net0.n_4_1_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_1_zneg.txt",net0.n_4_1_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_2_local.txt",net0.n_4_1_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_2_xpos.txt",net0.n_4_1_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_2_xneg.txt",net0.n_4_1_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_2_ypos.txt",net0.n_4_1_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_2_yneg.txt",net0.n_4_1_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_2_zpos.txt",net0.n_4_1_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_2_zneg.txt",net0.n_4_1_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_2_xpos.txt",net0.n_4_1_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_2_xneg.txt",net0.n_4_1_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_2_ypos.txt",net0.n_4_1_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_2_yneg.txt",net0.n_4_1_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_2_zpos.txt",net0.n_4_1_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_2_zneg.txt",net0.n_4_1_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_2_xpos.txt",net0.n_4_1_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_2_xneg.txt",net0.n_4_1_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_2_ypos.txt",net0.n_4_1_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_2_yneg.txt",net0.n_4_1_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_2_zpos.txt",net0.n_4_1_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_2_zneg.txt",net0.n_4_1_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_3_local.txt",net0.n_4_1_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_3_xpos.txt",net0.n_4_1_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_3_xneg.txt",net0.n_4_1_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_3_ypos.txt",net0.n_4_1_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_3_yneg.txt",net0.n_4_1_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_3_zpos.txt",net0.n_4_1_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_3_zneg.txt",net0.n_4_1_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_3_xpos.txt",net0.n_4_1_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_3_xneg.txt",net0.n_4_1_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_3_ypos.txt",net0.n_4_1_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_3_yneg.txt",net0.n_4_1_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_3_zpos.txt",net0.n_4_1_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_3_zneg.txt",net0.n_4_1_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_3_xpos.txt",net0.n_4_1_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_3_xneg.txt",net0.n_4_1_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_3_ypos.txt",net0.n_4_1_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_3_yneg.txt",net0.n_4_1_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_3_zpos.txt",net0.n_4_1_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_3_zneg.txt",net0.n_4_1_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_4_local.txt",net0.n_4_1_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_4_xpos.txt",net0.n_4_1_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_4_xneg.txt",net0.n_4_1_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_4_ypos.txt",net0.n_4_1_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_4_yneg.txt",net0.n_4_1_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_4_zpos.txt",net0.n_4_1_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_4_zneg.txt",net0.n_4_1_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_4_xpos.txt",net0.n_4_1_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_4_xneg.txt",net0.n_4_1_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_4_ypos.txt",net0.n_4_1_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_4_yneg.txt",net0.n_4_1_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_4_zpos.txt",net0.n_4_1_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_4_zneg.txt",net0.n_4_1_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_4_xpos.txt",net0.n_4_1_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_4_xneg.txt",net0.n_4_1_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_4_ypos.txt",net0.n_4_1_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_4_yneg.txt",net0.n_4_1_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_4_zpos.txt",net0.n_4_1_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_4_zneg.txt",net0.n_4_1_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_5_local.txt",net0.n_4_1_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_5_xpos.txt",net0.n_4_1_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_5_xneg.txt",net0.n_4_1_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_5_ypos.txt",net0.n_4_1_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_5_yneg.txt",net0.n_4_1_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_5_zpos.txt",net0.n_4_1_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_5_zneg.txt",net0.n_4_1_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_5_xpos.txt",net0.n_4_1_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_5_xneg.txt",net0.n_4_1_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_5_ypos.txt",net0.n_4_1_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_5_yneg.txt",net0.n_4_1_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_5_zpos.txt",net0.n_4_1_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_5_zneg.txt",net0.n_4_1_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_5_xpos.txt",net0.n_4_1_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_5_xneg.txt",net0.n_4_1_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_5_ypos.txt",net0.n_4_1_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_5_yneg.txt",net0.n_4_1_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_5_zpos.txt",net0.n_4_1_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_5_zneg.txt",net0.n_4_1_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_6_local.txt",net0.n_4_1_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_6_xpos.txt",net0.n_4_1_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_6_xneg.txt",net0.n_4_1_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_6_ypos.txt",net0.n_4_1_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_6_yneg.txt",net0.n_4_1_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_6_zpos.txt",net0.n_4_1_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_6_zneg.txt",net0.n_4_1_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_6_xpos.txt",net0.n_4_1_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_6_xneg.txt",net0.n_4_1_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_6_ypos.txt",net0.n_4_1_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_6_yneg.txt",net0.n_4_1_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_6_zpos.txt",net0.n_4_1_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_6_zneg.txt",net0.n_4_1_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_6_xpos.txt",net0.n_4_1_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_6_xneg.txt",net0.n_4_1_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_6_ypos.txt",net0.n_4_1_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_6_yneg.txt",net0.n_4_1_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_6_zpos.txt",net0.n_4_1_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_6_zneg.txt",net0.n_4_1_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_7_local.txt",net0.n_4_1_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_7_xpos.txt",net0.n_4_1_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_7_xneg.txt",net0.n_4_1_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_7_ypos.txt",net0.n_4_1_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_7_yneg.txt",net0.n_4_1_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_7_zpos.txt",net0.n_4_1_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_1_7_zneg.txt",net0.n_4_1_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_7_xpos.txt",net0.n_4_1_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_7_xneg.txt",net0.n_4_1_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_7_ypos.txt",net0.n_4_1_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_7_yneg.txt",net0.n_4_1_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_7_zpos.txt",net0.n_4_1_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_1_7_zneg.txt",net0.n_4_1_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_7_xpos.txt",net0.n_4_1_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_7_xneg.txt",net0.n_4_1_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_7_ypos.txt",net0.n_4_1_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_7_yneg.txt",net0.n_4_1_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_7_zpos.txt",net0.n_4_1_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_1_7_zneg.txt",net0.n_4_1_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_0_local.txt",net0.n_4_2_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_0_xpos.txt",net0.n_4_2_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_0_xneg.txt",net0.n_4_2_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_0_ypos.txt",net0.n_4_2_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_0_yneg.txt",net0.n_4_2_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_0_zpos.txt",net0.n_4_2_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_0_zneg.txt",net0.n_4_2_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_0_xpos.txt",net0.n_4_2_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_0_xneg.txt",net0.n_4_2_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_0_ypos.txt",net0.n_4_2_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_0_yneg.txt",net0.n_4_2_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_0_zpos.txt",net0.n_4_2_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_0_zneg.txt",net0.n_4_2_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_0_xpos.txt",net0.n_4_2_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_0_xneg.txt",net0.n_4_2_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_0_ypos.txt",net0.n_4_2_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_0_yneg.txt",net0.n_4_2_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_0_zpos.txt",net0.n_4_2_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_0_zneg.txt",net0.n_4_2_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_1_local.txt",net0.n_4_2_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_1_xpos.txt",net0.n_4_2_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_1_xneg.txt",net0.n_4_2_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_1_ypos.txt",net0.n_4_2_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_1_yneg.txt",net0.n_4_2_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_1_zpos.txt",net0.n_4_2_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_1_zneg.txt",net0.n_4_2_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_1_xpos.txt",net0.n_4_2_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_1_xneg.txt",net0.n_4_2_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_1_ypos.txt",net0.n_4_2_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_1_yneg.txt",net0.n_4_2_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_1_zpos.txt",net0.n_4_2_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_1_zneg.txt",net0.n_4_2_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_1_xpos.txt",net0.n_4_2_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_1_xneg.txt",net0.n_4_2_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_1_ypos.txt",net0.n_4_2_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_1_yneg.txt",net0.n_4_2_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_1_zpos.txt",net0.n_4_2_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_1_zneg.txt",net0.n_4_2_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_2_local.txt",net0.n_4_2_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_2_xpos.txt",net0.n_4_2_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_2_xneg.txt",net0.n_4_2_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_2_ypos.txt",net0.n_4_2_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_2_yneg.txt",net0.n_4_2_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_2_zpos.txt",net0.n_4_2_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_2_zneg.txt",net0.n_4_2_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_2_xpos.txt",net0.n_4_2_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_2_xneg.txt",net0.n_4_2_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_2_ypos.txt",net0.n_4_2_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_2_yneg.txt",net0.n_4_2_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_2_zpos.txt",net0.n_4_2_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_2_zneg.txt",net0.n_4_2_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_2_xpos.txt",net0.n_4_2_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_2_xneg.txt",net0.n_4_2_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_2_ypos.txt",net0.n_4_2_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_2_yneg.txt",net0.n_4_2_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_2_zpos.txt",net0.n_4_2_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_2_zneg.txt",net0.n_4_2_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_3_local.txt",net0.n_4_2_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_3_xpos.txt",net0.n_4_2_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_3_xneg.txt",net0.n_4_2_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_3_ypos.txt",net0.n_4_2_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_3_yneg.txt",net0.n_4_2_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_3_zpos.txt",net0.n_4_2_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_3_zneg.txt",net0.n_4_2_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_3_xpos.txt",net0.n_4_2_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_3_xneg.txt",net0.n_4_2_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_3_ypos.txt",net0.n_4_2_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_3_yneg.txt",net0.n_4_2_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_3_zpos.txt",net0.n_4_2_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_3_zneg.txt",net0.n_4_2_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_3_xpos.txt",net0.n_4_2_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_3_xneg.txt",net0.n_4_2_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_3_ypos.txt",net0.n_4_2_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_3_yneg.txt",net0.n_4_2_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_3_zpos.txt",net0.n_4_2_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_3_zneg.txt",net0.n_4_2_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_4_local.txt",net0.n_4_2_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_4_xpos.txt",net0.n_4_2_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_4_xneg.txt",net0.n_4_2_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_4_ypos.txt",net0.n_4_2_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_4_yneg.txt",net0.n_4_2_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_4_zpos.txt",net0.n_4_2_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_4_zneg.txt",net0.n_4_2_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_4_xpos.txt",net0.n_4_2_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_4_xneg.txt",net0.n_4_2_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_4_ypos.txt",net0.n_4_2_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_4_yneg.txt",net0.n_4_2_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_4_zpos.txt",net0.n_4_2_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_4_zneg.txt",net0.n_4_2_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_4_xpos.txt",net0.n_4_2_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_4_xneg.txt",net0.n_4_2_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_4_ypos.txt",net0.n_4_2_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_4_yneg.txt",net0.n_4_2_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_4_zpos.txt",net0.n_4_2_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_4_zneg.txt",net0.n_4_2_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_5_local.txt",net0.n_4_2_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_5_xpos.txt",net0.n_4_2_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_5_xneg.txt",net0.n_4_2_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_5_ypos.txt",net0.n_4_2_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_5_yneg.txt",net0.n_4_2_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_5_zpos.txt",net0.n_4_2_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_5_zneg.txt",net0.n_4_2_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_5_xpos.txt",net0.n_4_2_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_5_xneg.txt",net0.n_4_2_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_5_ypos.txt",net0.n_4_2_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_5_yneg.txt",net0.n_4_2_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_5_zpos.txt",net0.n_4_2_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_5_zneg.txt",net0.n_4_2_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_5_xpos.txt",net0.n_4_2_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_5_xneg.txt",net0.n_4_2_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_5_ypos.txt",net0.n_4_2_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_5_yneg.txt",net0.n_4_2_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_5_zpos.txt",net0.n_4_2_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_5_zneg.txt",net0.n_4_2_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_6_local.txt",net0.n_4_2_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_6_xpos.txt",net0.n_4_2_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_6_xneg.txt",net0.n_4_2_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_6_ypos.txt",net0.n_4_2_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_6_yneg.txt",net0.n_4_2_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_6_zpos.txt",net0.n_4_2_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_6_zneg.txt",net0.n_4_2_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_6_xpos.txt",net0.n_4_2_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_6_xneg.txt",net0.n_4_2_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_6_ypos.txt",net0.n_4_2_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_6_yneg.txt",net0.n_4_2_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_6_zpos.txt",net0.n_4_2_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_6_zneg.txt",net0.n_4_2_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_6_xpos.txt",net0.n_4_2_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_6_xneg.txt",net0.n_4_2_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_6_ypos.txt",net0.n_4_2_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_6_yneg.txt",net0.n_4_2_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_6_zpos.txt",net0.n_4_2_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_6_zneg.txt",net0.n_4_2_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_7_local.txt",net0.n_4_2_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_7_xpos.txt",net0.n_4_2_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_7_xneg.txt",net0.n_4_2_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_7_ypos.txt",net0.n_4_2_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_7_yneg.txt",net0.n_4_2_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_7_zpos.txt",net0.n_4_2_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_2_7_zneg.txt",net0.n_4_2_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_7_xpos.txt",net0.n_4_2_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_7_xneg.txt",net0.n_4_2_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_7_ypos.txt",net0.n_4_2_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_7_yneg.txt",net0.n_4_2_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_7_zpos.txt",net0.n_4_2_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_2_7_zneg.txt",net0.n_4_2_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_7_xpos.txt",net0.n_4_2_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_7_xneg.txt",net0.n_4_2_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_7_ypos.txt",net0.n_4_2_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_7_yneg.txt",net0.n_4_2_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_7_zpos.txt",net0.n_4_2_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_2_7_zneg.txt",net0.n_4_2_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_0_local.txt",net0.n_4_3_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_0_xpos.txt",net0.n_4_3_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_0_xneg.txt",net0.n_4_3_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_0_ypos.txt",net0.n_4_3_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_0_yneg.txt",net0.n_4_3_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_0_zpos.txt",net0.n_4_3_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_0_zneg.txt",net0.n_4_3_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_0_xpos.txt",net0.n_4_3_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_0_xneg.txt",net0.n_4_3_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_0_ypos.txt",net0.n_4_3_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_0_yneg.txt",net0.n_4_3_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_0_zpos.txt",net0.n_4_3_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_0_zneg.txt",net0.n_4_3_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_0_xpos.txt",net0.n_4_3_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_0_xneg.txt",net0.n_4_3_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_0_ypos.txt",net0.n_4_3_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_0_yneg.txt",net0.n_4_3_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_0_zpos.txt",net0.n_4_3_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_0_zneg.txt",net0.n_4_3_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_1_local.txt",net0.n_4_3_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_1_xpos.txt",net0.n_4_3_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_1_xneg.txt",net0.n_4_3_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_1_ypos.txt",net0.n_4_3_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_1_yneg.txt",net0.n_4_3_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_1_zpos.txt",net0.n_4_3_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_1_zneg.txt",net0.n_4_3_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_1_xpos.txt",net0.n_4_3_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_1_xneg.txt",net0.n_4_3_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_1_ypos.txt",net0.n_4_3_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_1_yneg.txt",net0.n_4_3_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_1_zpos.txt",net0.n_4_3_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_1_zneg.txt",net0.n_4_3_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_1_xpos.txt",net0.n_4_3_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_1_xneg.txt",net0.n_4_3_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_1_ypos.txt",net0.n_4_3_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_1_yneg.txt",net0.n_4_3_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_1_zpos.txt",net0.n_4_3_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_1_zneg.txt",net0.n_4_3_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_2_local.txt",net0.n_4_3_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_2_xpos.txt",net0.n_4_3_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_2_xneg.txt",net0.n_4_3_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_2_ypos.txt",net0.n_4_3_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_2_yneg.txt",net0.n_4_3_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_2_zpos.txt",net0.n_4_3_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_2_zneg.txt",net0.n_4_3_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_2_xpos.txt",net0.n_4_3_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_2_xneg.txt",net0.n_4_3_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_2_ypos.txt",net0.n_4_3_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_2_yneg.txt",net0.n_4_3_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_2_zpos.txt",net0.n_4_3_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_2_zneg.txt",net0.n_4_3_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_2_xpos.txt",net0.n_4_3_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_2_xneg.txt",net0.n_4_3_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_2_ypos.txt",net0.n_4_3_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_2_yneg.txt",net0.n_4_3_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_2_zpos.txt",net0.n_4_3_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_2_zneg.txt",net0.n_4_3_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_3_local.txt",net0.n_4_3_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_3_xpos.txt",net0.n_4_3_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_3_xneg.txt",net0.n_4_3_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_3_ypos.txt",net0.n_4_3_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_3_yneg.txt",net0.n_4_3_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_3_zpos.txt",net0.n_4_3_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_3_zneg.txt",net0.n_4_3_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_3_xpos.txt",net0.n_4_3_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_3_xneg.txt",net0.n_4_3_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_3_ypos.txt",net0.n_4_3_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_3_yneg.txt",net0.n_4_3_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_3_zpos.txt",net0.n_4_3_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_3_zneg.txt",net0.n_4_3_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_3_xpos.txt",net0.n_4_3_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_3_xneg.txt",net0.n_4_3_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_3_ypos.txt",net0.n_4_3_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_3_yneg.txt",net0.n_4_3_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_3_zpos.txt",net0.n_4_3_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_3_zneg.txt",net0.n_4_3_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_4_local.txt",net0.n_4_3_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_4_xpos.txt",net0.n_4_3_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_4_xneg.txt",net0.n_4_3_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_4_ypos.txt",net0.n_4_3_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_4_yneg.txt",net0.n_4_3_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_4_zpos.txt",net0.n_4_3_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_4_zneg.txt",net0.n_4_3_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_4_xpos.txt",net0.n_4_3_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_4_xneg.txt",net0.n_4_3_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_4_ypos.txt",net0.n_4_3_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_4_yneg.txt",net0.n_4_3_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_4_zpos.txt",net0.n_4_3_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_4_zneg.txt",net0.n_4_3_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_4_xpos.txt",net0.n_4_3_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_4_xneg.txt",net0.n_4_3_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_4_ypos.txt",net0.n_4_3_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_4_yneg.txt",net0.n_4_3_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_4_zpos.txt",net0.n_4_3_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_4_zneg.txt",net0.n_4_3_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_5_local.txt",net0.n_4_3_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_5_xpos.txt",net0.n_4_3_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_5_xneg.txt",net0.n_4_3_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_5_ypos.txt",net0.n_4_3_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_5_yneg.txt",net0.n_4_3_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_5_zpos.txt",net0.n_4_3_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_5_zneg.txt",net0.n_4_3_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_5_xpos.txt",net0.n_4_3_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_5_xneg.txt",net0.n_4_3_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_5_ypos.txt",net0.n_4_3_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_5_yneg.txt",net0.n_4_3_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_5_zpos.txt",net0.n_4_3_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_5_zneg.txt",net0.n_4_3_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_5_xpos.txt",net0.n_4_3_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_5_xneg.txt",net0.n_4_3_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_5_ypos.txt",net0.n_4_3_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_5_yneg.txt",net0.n_4_3_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_5_zpos.txt",net0.n_4_3_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_5_zneg.txt",net0.n_4_3_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_6_local.txt",net0.n_4_3_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_6_xpos.txt",net0.n_4_3_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_6_xneg.txt",net0.n_4_3_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_6_ypos.txt",net0.n_4_3_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_6_yneg.txt",net0.n_4_3_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_6_zpos.txt",net0.n_4_3_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_6_zneg.txt",net0.n_4_3_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_6_xpos.txt",net0.n_4_3_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_6_xneg.txt",net0.n_4_3_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_6_ypos.txt",net0.n_4_3_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_6_yneg.txt",net0.n_4_3_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_6_zpos.txt",net0.n_4_3_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_6_zneg.txt",net0.n_4_3_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_6_xpos.txt",net0.n_4_3_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_6_xneg.txt",net0.n_4_3_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_6_ypos.txt",net0.n_4_3_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_6_yneg.txt",net0.n_4_3_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_6_zpos.txt",net0.n_4_3_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_6_zneg.txt",net0.n_4_3_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_7_local.txt",net0.n_4_3_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_7_xpos.txt",net0.n_4_3_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_7_xneg.txt",net0.n_4_3_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_7_ypos.txt",net0.n_4_3_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_7_yneg.txt",net0.n_4_3_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_7_zpos.txt",net0.n_4_3_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_3_7_zneg.txt",net0.n_4_3_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_7_xpos.txt",net0.n_4_3_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_7_xneg.txt",net0.n_4_3_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_7_ypos.txt",net0.n_4_3_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_7_yneg.txt",net0.n_4_3_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_7_zpos.txt",net0.n_4_3_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_3_7_zneg.txt",net0.n_4_3_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_7_xpos.txt",net0.n_4_3_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_7_xneg.txt",net0.n_4_3_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_7_ypos.txt",net0.n_4_3_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_7_yneg.txt",net0.n_4_3_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_7_zpos.txt",net0.n_4_3_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_3_7_zneg.txt",net0.n_4_3_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_0_local.txt",net0.n_4_4_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_0_xpos.txt",net0.n_4_4_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_0_xneg.txt",net0.n_4_4_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_0_ypos.txt",net0.n_4_4_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_0_yneg.txt",net0.n_4_4_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_0_zpos.txt",net0.n_4_4_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_0_zneg.txt",net0.n_4_4_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_0_xpos.txt",net0.n_4_4_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_0_xneg.txt",net0.n_4_4_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_0_ypos.txt",net0.n_4_4_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_0_yneg.txt",net0.n_4_4_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_0_zpos.txt",net0.n_4_4_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_0_zneg.txt",net0.n_4_4_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_0_xpos.txt",net0.n_4_4_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_0_xneg.txt",net0.n_4_4_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_0_ypos.txt",net0.n_4_4_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_0_yneg.txt",net0.n_4_4_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_0_zpos.txt",net0.n_4_4_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_0_zneg.txt",net0.n_4_4_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_1_local.txt",net0.n_4_4_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_1_xpos.txt",net0.n_4_4_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_1_xneg.txt",net0.n_4_4_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_1_ypos.txt",net0.n_4_4_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_1_yneg.txt",net0.n_4_4_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_1_zpos.txt",net0.n_4_4_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_1_zneg.txt",net0.n_4_4_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_1_xpos.txt",net0.n_4_4_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_1_xneg.txt",net0.n_4_4_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_1_ypos.txt",net0.n_4_4_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_1_yneg.txt",net0.n_4_4_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_1_zpos.txt",net0.n_4_4_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_1_zneg.txt",net0.n_4_4_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_1_xpos.txt",net0.n_4_4_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_1_xneg.txt",net0.n_4_4_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_1_ypos.txt",net0.n_4_4_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_1_yneg.txt",net0.n_4_4_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_1_zpos.txt",net0.n_4_4_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_1_zneg.txt",net0.n_4_4_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_2_local.txt",net0.n_4_4_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_2_xpos.txt",net0.n_4_4_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_2_xneg.txt",net0.n_4_4_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_2_ypos.txt",net0.n_4_4_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_2_yneg.txt",net0.n_4_4_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_2_zpos.txt",net0.n_4_4_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_2_zneg.txt",net0.n_4_4_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_2_xpos.txt",net0.n_4_4_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_2_xneg.txt",net0.n_4_4_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_2_ypos.txt",net0.n_4_4_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_2_yneg.txt",net0.n_4_4_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_2_zpos.txt",net0.n_4_4_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_2_zneg.txt",net0.n_4_4_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_2_xpos.txt",net0.n_4_4_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_2_xneg.txt",net0.n_4_4_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_2_ypos.txt",net0.n_4_4_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_2_yneg.txt",net0.n_4_4_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_2_zpos.txt",net0.n_4_4_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_2_zneg.txt",net0.n_4_4_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_3_local.txt",net0.n_4_4_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_3_xpos.txt",net0.n_4_4_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_3_xneg.txt",net0.n_4_4_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_3_ypos.txt",net0.n_4_4_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_3_yneg.txt",net0.n_4_4_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_3_zpos.txt",net0.n_4_4_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_3_zneg.txt",net0.n_4_4_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_3_xpos.txt",net0.n_4_4_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_3_xneg.txt",net0.n_4_4_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_3_ypos.txt",net0.n_4_4_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_3_yneg.txt",net0.n_4_4_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_3_zpos.txt",net0.n_4_4_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_3_zneg.txt",net0.n_4_4_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_3_xpos.txt",net0.n_4_4_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_3_xneg.txt",net0.n_4_4_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_3_ypos.txt",net0.n_4_4_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_3_yneg.txt",net0.n_4_4_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_3_zpos.txt",net0.n_4_4_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_3_zneg.txt",net0.n_4_4_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_4_local.txt",net0.n_4_4_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_4_xpos.txt",net0.n_4_4_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_4_xneg.txt",net0.n_4_4_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_4_ypos.txt",net0.n_4_4_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_4_yneg.txt",net0.n_4_4_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_4_zpos.txt",net0.n_4_4_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_4_zneg.txt",net0.n_4_4_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_4_xpos.txt",net0.n_4_4_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_4_xneg.txt",net0.n_4_4_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_4_ypos.txt",net0.n_4_4_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_4_yneg.txt",net0.n_4_4_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_4_zpos.txt",net0.n_4_4_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_4_zneg.txt",net0.n_4_4_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_4_xpos.txt",net0.n_4_4_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_4_xneg.txt",net0.n_4_4_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_4_ypos.txt",net0.n_4_4_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_4_yneg.txt",net0.n_4_4_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_4_zpos.txt",net0.n_4_4_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_4_zneg.txt",net0.n_4_4_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_5_local.txt",net0.n_4_4_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_5_xpos.txt",net0.n_4_4_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_5_xneg.txt",net0.n_4_4_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_5_ypos.txt",net0.n_4_4_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_5_yneg.txt",net0.n_4_4_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_5_zpos.txt",net0.n_4_4_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_5_zneg.txt",net0.n_4_4_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_5_xpos.txt",net0.n_4_4_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_5_xneg.txt",net0.n_4_4_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_5_ypos.txt",net0.n_4_4_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_5_yneg.txt",net0.n_4_4_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_5_zpos.txt",net0.n_4_4_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_5_zneg.txt",net0.n_4_4_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_5_xpos.txt",net0.n_4_4_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_5_xneg.txt",net0.n_4_4_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_5_ypos.txt",net0.n_4_4_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_5_yneg.txt",net0.n_4_4_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_5_zpos.txt",net0.n_4_4_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_5_zneg.txt",net0.n_4_4_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_6_local.txt",net0.n_4_4_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_6_xpos.txt",net0.n_4_4_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_6_xneg.txt",net0.n_4_4_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_6_ypos.txt",net0.n_4_4_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_6_yneg.txt",net0.n_4_4_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_6_zpos.txt",net0.n_4_4_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_6_zneg.txt",net0.n_4_4_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_6_xpos.txt",net0.n_4_4_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_6_xneg.txt",net0.n_4_4_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_6_ypos.txt",net0.n_4_4_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_6_yneg.txt",net0.n_4_4_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_6_zpos.txt",net0.n_4_4_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_6_zneg.txt",net0.n_4_4_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_6_xpos.txt",net0.n_4_4_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_6_xneg.txt",net0.n_4_4_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_6_ypos.txt",net0.n_4_4_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_6_yneg.txt",net0.n_4_4_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_6_zpos.txt",net0.n_4_4_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_6_zneg.txt",net0.n_4_4_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_7_local.txt",net0.n_4_4_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_7_xpos.txt",net0.n_4_4_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_7_xneg.txt",net0.n_4_4_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_7_ypos.txt",net0.n_4_4_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_7_yneg.txt",net0.n_4_4_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_7_zpos.txt",net0.n_4_4_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_4_7_zneg.txt",net0.n_4_4_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_7_xpos.txt",net0.n_4_4_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_7_xneg.txt",net0.n_4_4_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_7_ypos.txt",net0.n_4_4_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_7_yneg.txt",net0.n_4_4_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_7_zpos.txt",net0.n_4_4_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_4_7_zneg.txt",net0.n_4_4_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_7_xpos.txt",net0.n_4_4_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_7_xneg.txt",net0.n_4_4_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_7_ypos.txt",net0.n_4_4_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_7_yneg.txt",net0.n_4_4_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_7_zpos.txt",net0.n_4_4_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_4_7_zneg.txt",net0.n_4_4_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_0_local.txt",net0.n_4_5_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_0_xpos.txt",net0.n_4_5_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_0_xneg.txt",net0.n_4_5_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_0_ypos.txt",net0.n_4_5_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_0_yneg.txt",net0.n_4_5_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_0_zpos.txt",net0.n_4_5_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_0_zneg.txt",net0.n_4_5_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_0_xpos.txt",net0.n_4_5_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_0_xneg.txt",net0.n_4_5_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_0_ypos.txt",net0.n_4_5_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_0_yneg.txt",net0.n_4_5_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_0_zpos.txt",net0.n_4_5_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_0_zneg.txt",net0.n_4_5_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_0_xpos.txt",net0.n_4_5_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_0_xneg.txt",net0.n_4_5_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_0_ypos.txt",net0.n_4_5_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_0_yneg.txt",net0.n_4_5_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_0_zpos.txt",net0.n_4_5_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_0_zneg.txt",net0.n_4_5_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_1_local.txt",net0.n_4_5_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_1_xpos.txt",net0.n_4_5_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_1_xneg.txt",net0.n_4_5_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_1_ypos.txt",net0.n_4_5_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_1_yneg.txt",net0.n_4_5_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_1_zpos.txt",net0.n_4_5_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_1_zneg.txt",net0.n_4_5_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_1_xpos.txt",net0.n_4_5_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_1_xneg.txt",net0.n_4_5_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_1_ypos.txt",net0.n_4_5_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_1_yneg.txt",net0.n_4_5_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_1_zpos.txt",net0.n_4_5_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_1_zneg.txt",net0.n_4_5_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_1_xpos.txt",net0.n_4_5_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_1_xneg.txt",net0.n_4_5_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_1_ypos.txt",net0.n_4_5_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_1_yneg.txt",net0.n_4_5_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_1_zpos.txt",net0.n_4_5_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_1_zneg.txt",net0.n_4_5_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_2_local.txt",net0.n_4_5_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_2_xpos.txt",net0.n_4_5_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_2_xneg.txt",net0.n_4_5_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_2_ypos.txt",net0.n_4_5_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_2_yneg.txt",net0.n_4_5_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_2_zpos.txt",net0.n_4_5_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_2_zneg.txt",net0.n_4_5_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_2_xpos.txt",net0.n_4_5_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_2_xneg.txt",net0.n_4_5_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_2_ypos.txt",net0.n_4_5_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_2_yneg.txt",net0.n_4_5_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_2_zpos.txt",net0.n_4_5_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_2_zneg.txt",net0.n_4_5_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_2_xpos.txt",net0.n_4_5_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_2_xneg.txt",net0.n_4_5_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_2_ypos.txt",net0.n_4_5_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_2_yneg.txt",net0.n_4_5_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_2_zpos.txt",net0.n_4_5_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_2_zneg.txt",net0.n_4_5_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_3_local.txt",net0.n_4_5_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_3_xpos.txt",net0.n_4_5_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_3_xneg.txt",net0.n_4_5_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_3_ypos.txt",net0.n_4_5_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_3_yneg.txt",net0.n_4_5_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_3_zpos.txt",net0.n_4_5_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_3_zneg.txt",net0.n_4_5_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_3_xpos.txt",net0.n_4_5_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_3_xneg.txt",net0.n_4_5_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_3_ypos.txt",net0.n_4_5_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_3_yneg.txt",net0.n_4_5_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_3_zpos.txt",net0.n_4_5_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_3_zneg.txt",net0.n_4_5_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_3_xpos.txt",net0.n_4_5_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_3_xneg.txt",net0.n_4_5_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_3_ypos.txt",net0.n_4_5_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_3_yneg.txt",net0.n_4_5_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_3_zpos.txt",net0.n_4_5_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_3_zneg.txt",net0.n_4_5_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_4_local.txt",net0.n_4_5_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_4_xpos.txt",net0.n_4_5_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_4_xneg.txt",net0.n_4_5_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_4_ypos.txt",net0.n_4_5_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_4_yneg.txt",net0.n_4_5_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_4_zpos.txt",net0.n_4_5_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_4_zneg.txt",net0.n_4_5_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_4_xpos.txt",net0.n_4_5_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_4_xneg.txt",net0.n_4_5_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_4_ypos.txt",net0.n_4_5_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_4_yneg.txt",net0.n_4_5_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_4_zpos.txt",net0.n_4_5_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_4_zneg.txt",net0.n_4_5_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_4_xpos.txt",net0.n_4_5_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_4_xneg.txt",net0.n_4_5_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_4_ypos.txt",net0.n_4_5_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_4_yneg.txt",net0.n_4_5_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_4_zpos.txt",net0.n_4_5_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_4_zneg.txt",net0.n_4_5_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_5_local.txt",net0.n_4_5_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_5_xpos.txt",net0.n_4_5_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_5_xneg.txt",net0.n_4_5_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_5_ypos.txt",net0.n_4_5_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_5_yneg.txt",net0.n_4_5_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_5_zpos.txt",net0.n_4_5_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_5_zneg.txt",net0.n_4_5_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_5_xpos.txt",net0.n_4_5_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_5_xneg.txt",net0.n_4_5_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_5_ypos.txt",net0.n_4_5_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_5_yneg.txt",net0.n_4_5_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_5_zpos.txt",net0.n_4_5_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_5_zneg.txt",net0.n_4_5_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_5_xpos.txt",net0.n_4_5_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_5_xneg.txt",net0.n_4_5_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_5_ypos.txt",net0.n_4_5_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_5_yneg.txt",net0.n_4_5_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_5_zpos.txt",net0.n_4_5_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_5_zneg.txt",net0.n_4_5_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_6_local.txt",net0.n_4_5_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_6_xpos.txt",net0.n_4_5_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_6_xneg.txt",net0.n_4_5_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_6_ypos.txt",net0.n_4_5_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_6_yneg.txt",net0.n_4_5_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_6_zpos.txt",net0.n_4_5_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_6_zneg.txt",net0.n_4_5_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_6_xpos.txt",net0.n_4_5_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_6_xneg.txt",net0.n_4_5_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_6_ypos.txt",net0.n_4_5_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_6_yneg.txt",net0.n_4_5_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_6_zpos.txt",net0.n_4_5_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_6_zneg.txt",net0.n_4_5_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_6_xpos.txt",net0.n_4_5_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_6_xneg.txt",net0.n_4_5_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_6_ypos.txt",net0.n_4_5_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_6_yneg.txt",net0.n_4_5_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_6_zpos.txt",net0.n_4_5_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_6_zneg.txt",net0.n_4_5_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_7_local.txt",net0.n_4_5_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_7_xpos.txt",net0.n_4_5_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_7_xneg.txt",net0.n_4_5_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_7_ypos.txt",net0.n_4_5_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_7_yneg.txt",net0.n_4_5_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_7_zpos.txt",net0.n_4_5_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_5_7_zneg.txt",net0.n_4_5_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_7_xpos.txt",net0.n_4_5_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_7_xneg.txt",net0.n_4_5_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_7_ypos.txt",net0.n_4_5_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_7_yneg.txt",net0.n_4_5_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_7_zpos.txt",net0.n_4_5_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_5_7_zneg.txt",net0.n_4_5_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_7_xpos.txt",net0.n_4_5_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_7_xneg.txt",net0.n_4_5_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_7_ypos.txt",net0.n_4_5_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_7_yneg.txt",net0.n_4_5_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_7_zpos.txt",net0.n_4_5_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_5_7_zneg.txt",net0.n_4_5_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_0_local.txt",net0.n_4_6_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_0_xpos.txt",net0.n_4_6_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_0_xneg.txt",net0.n_4_6_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_0_ypos.txt",net0.n_4_6_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_0_yneg.txt",net0.n_4_6_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_0_zpos.txt",net0.n_4_6_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_0_zneg.txt",net0.n_4_6_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_0_xpos.txt",net0.n_4_6_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_0_xneg.txt",net0.n_4_6_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_0_ypos.txt",net0.n_4_6_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_0_yneg.txt",net0.n_4_6_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_0_zpos.txt",net0.n_4_6_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_0_zneg.txt",net0.n_4_6_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_0_xpos.txt",net0.n_4_6_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_0_xneg.txt",net0.n_4_6_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_0_ypos.txt",net0.n_4_6_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_0_yneg.txt",net0.n_4_6_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_0_zpos.txt",net0.n_4_6_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_0_zneg.txt",net0.n_4_6_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_1_local.txt",net0.n_4_6_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_1_xpos.txt",net0.n_4_6_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_1_xneg.txt",net0.n_4_6_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_1_ypos.txt",net0.n_4_6_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_1_yneg.txt",net0.n_4_6_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_1_zpos.txt",net0.n_4_6_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_1_zneg.txt",net0.n_4_6_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_1_xpos.txt",net0.n_4_6_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_1_xneg.txt",net0.n_4_6_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_1_ypos.txt",net0.n_4_6_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_1_yneg.txt",net0.n_4_6_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_1_zpos.txt",net0.n_4_6_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_1_zneg.txt",net0.n_4_6_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_1_xpos.txt",net0.n_4_6_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_1_xneg.txt",net0.n_4_6_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_1_ypos.txt",net0.n_4_6_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_1_yneg.txt",net0.n_4_6_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_1_zpos.txt",net0.n_4_6_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_1_zneg.txt",net0.n_4_6_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_2_local.txt",net0.n_4_6_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_2_xpos.txt",net0.n_4_6_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_2_xneg.txt",net0.n_4_6_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_2_ypos.txt",net0.n_4_6_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_2_yneg.txt",net0.n_4_6_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_2_zpos.txt",net0.n_4_6_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_2_zneg.txt",net0.n_4_6_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_2_xpos.txt",net0.n_4_6_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_2_xneg.txt",net0.n_4_6_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_2_ypos.txt",net0.n_4_6_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_2_yneg.txt",net0.n_4_6_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_2_zpos.txt",net0.n_4_6_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_2_zneg.txt",net0.n_4_6_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_2_xpos.txt",net0.n_4_6_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_2_xneg.txt",net0.n_4_6_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_2_ypos.txt",net0.n_4_6_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_2_yneg.txt",net0.n_4_6_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_2_zpos.txt",net0.n_4_6_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_2_zneg.txt",net0.n_4_6_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_3_local.txt",net0.n_4_6_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_3_xpos.txt",net0.n_4_6_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_3_xneg.txt",net0.n_4_6_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_3_ypos.txt",net0.n_4_6_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_3_yneg.txt",net0.n_4_6_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_3_zpos.txt",net0.n_4_6_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_3_zneg.txt",net0.n_4_6_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_3_xpos.txt",net0.n_4_6_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_3_xneg.txt",net0.n_4_6_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_3_ypos.txt",net0.n_4_6_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_3_yneg.txt",net0.n_4_6_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_3_zpos.txt",net0.n_4_6_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_3_zneg.txt",net0.n_4_6_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_3_xpos.txt",net0.n_4_6_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_3_xneg.txt",net0.n_4_6_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_3_ypos.txt",net0.n_4_6_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_3_yneg.txt",net0.n_4_6_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_3_zpos.txt",net0.n_4_6_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_3_zneg.txt",net0.n_4_6_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_4_local.txt",net0.n_4_6_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_4_xpos.txt",net0.n_4_6_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_4_xneg.txt",net0.n_4_6_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_4_ypos.txt",net0.n_4_6_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_4_yneg.txt",net0.n_4_6_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_4_zpos.txt",net0.n_4_6_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_4_zneg.txt",net0.n_4_6_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_4_xpos.txt",net0.n_4_6_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_4_xneg.txt",net0.n_4_6_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_4_ypos.txt",net0.n_4_6_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_4_yneg.txt",net0.n_4_6_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_4_zpos.txt",net0.n_4_6_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_4_zneg.txt",net0.n_4_6_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_4_xpos.txt",net0.n_4_6_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_4_xneg.txt",net0.n_4_6_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_4_ypos.txt",net0.n_4_6_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_4_yneg.txt",net0.n_4_6_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_4_zpos.txt",net0.n_4_6_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_4_zneg.txt",net0.n_4_6_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_5_local.txt",net0.n_4_6_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_5_xpos.txt",net0.n_4_6_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_5_xneg.txt",net0.n_4_6_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_5_ypos.txt",net0.n_4_6_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_5_yneg.txt",net0.n_4_6_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_5_zpos.txt",net0.n_4_6_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_5_zneg.txt",net0.n_4_6_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_5_xpos.txt",net0.n_4_6_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_5_xneg.txt",net0.n_4_6_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_5_ypos.txt",net0.n_4_6_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_5_yneg.txt",net0.n_4_6_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_5_zpos.txt",net0.n_4_6_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_5_zneg.txt",net0.n_4_6_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_5_xpos.txt",net0.n_4_6_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_5_xneg.txt",net0.n_4_6_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_5_ypos.txt",net0.n_4_6_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_5_yneg.txt",net0.n_4_6_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_5_zpos.txt",net0.n_4_6_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_5_zneg.txt",net0.n_4_6_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_6_local.txt",net0.n_4_6_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_6_xpos.txt",net0.n_4_6_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_6_xneg.txt",net0.n_4_6_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_6_ypos.txt",net0.n_4_6_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_6_yneg.txt",net0.n_4_6_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_6_zpos.txt",net0.n_4_6_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_6_zneg.txt",net0.n_4_6_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_6_xpos.txt",net0.n_4_6_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_6_xneg.txt",net0.n_4_6_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_6_ypos.txt",net0.n_4_6_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_6_yneg.txt",net0.n_4_6_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_6_zpos.txt",net0.n_4_6_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_6_zneg.txt",net0.n_4_6_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_6_xpos.txt",net0.n_4_6_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_6_xneg.txt",net0.n_4_6_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_6_ypos.txt",net0.n_4_6_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_6_yneg.txt",net0.n_4_6_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_6_zpos.txt",net0.n_4_6_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_6_zneg.txt",net0.n_4_6_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_7_local.txt",net0.n_4_6_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_7_xpos.txt",net0.n_4_6_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_7_xneg.txt",net0.n_4_6_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_7_ypos.txt",net0.n_4_6_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_7_yneg.txt",net0.n_4_6_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_7_zpos.txt",net0.n_4_6_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_6_7_zneg.txt",net0.n_4_6_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_7_xpos.txt",net0.n_4_6_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_7_xneg.txt",net0.n_4_6_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_7_ypos.txt",net0.n_4_6_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_7_yneg.txt",net0.n_4_6_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_7_zpos.txt",net0.n_4_6_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_6_7_zneg.txt",net0.n_4_6_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_7_xpos.txt",net0.n_4_6_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_7_xneg.txt",net0.n_4_6_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_7_ypos.txt",net0.n_4_6_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_7_yneg.txt",net0.n_4_6_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_7_zpos.txt",net0.n_4_6_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_6_7_zneg.txt",net0.n_4_6_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_0_local.txt",net0.n_4_7_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_0_xpos.txt",net0.n_4_7_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_0_xneg.txt",net0.n_4_7_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_0_ypos.txt",net0.n_4_7_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_0_yneg.txt",net0.n_4_7_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_0_zpos.txt",net0.n_4_7_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_0_zneg.txt",net0.n_4_7_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_0_xpos.txt",net0.n_4_7_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_0_xneg.txt",net0.n_4_7_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_0_ypos.txt",net0.n_4_7_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_0_yneg.txt",net0.n_4_7_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_0_zpos.txt",net0.n_4_7_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_0_zneg.txt",net0.n_4_7_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_0_xpos.txt",net0.n_4_7_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_0_xneg.txt",net0.n_4_7_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_0_ypos.txt",net0.n_4_7_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_0_yneg.txt",net0.n_4_7_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_0_zpos.txt",net0.n_4_7_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_0_zneg.txt",net0.n_4_7_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_1_local.txt",net0.n_4_7_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_1_xpos.txt",net0.n_4_7_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_1_xneg.txt",net0.n_4_7_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_1_ypos.txt",net0.n_4_7_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_1_yneg.txt",net0.n_4_7_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_1_zpos.txt",net0.n_4_7_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_1_zneg.txt",net0.n_4_7_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_1_xpos.txt",net0.n_4_7_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_1_xneg.txt",net0.n_4_7_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_1_ypos.txt",net0.n_4_7_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_1_yneg.txt",net0.n_4_7_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_1_zpos.txt",net0.n_4_7_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_1_zneg.txt",net0.n_4_7_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_1_xpos.txt",net0.n_4_7_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_1_xneg.txt",net0.n_4_7_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_1_ypos.txt",net0.n_4_7_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_1_yneg.txt",net0.n_4_7_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_1_zpos.txt",net0.n_4_7_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_1_zneg.txt",net0.n_4_7_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_2_local.txt",net0.n_4_7_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_2_xpos.txt",net0.n_4_7_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_2_xneg.txt",net0.n_4_7_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_2_ypos.txt",net0.n_4_7_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_2_yneg.txt",net0.n_4_7_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_2_zpos.txt",net0.n_4_7_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_2_zneg.txt",net0.n_4_7_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_2_xpos.txt",net0.n_4_7_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_2_xneg.txt",net0.n_4_7_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_2_ypos.txt",net0.n_4_7_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_2_yneg.txt",net0.n_4_7_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_2_zpos.txt",net0.n_4_7_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_2_zneg.txt",net0.n_4_7_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_2_xpos.txt",net0.n_4_7_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_2_xneg.txt",net0.n_4_7_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_2_ypos.txt",net0.n_4_7_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_2_yneg.txt",net0.n_4_7_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_2_zpos.txt",net0.n_4_7_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_2_zneg.txt",net0.n_4_7_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_3_local.txt",net0.n_4_7_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_3_xpos.txt",net0.n_4_7_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_3_xneg.txt",net0.n_4_7_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_3_ypos.txt",net0.n_4_7_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_3_yneg.txt",net0.n_4_7_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_3_zpos.txt",net0.n_4_7_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_3_zneg.txt",net0.n_4_7_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_3_xpos.txt",net0.n_4_7_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_3_xneg.txt",net0.n_4_7_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_3_ypos.txt",net0.n_4_7_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_3_yneg.txt",net0.n_4_7_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_3_zpos.txt",net0.n_4_7_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_3_zneg.txt",net0.n_4_7_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_3_xpos.txt",net0.n_4_7_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_3_xneg.txt",net0.n_4_7_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_3_ypos.txt",net0.n_4_7_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_3_yneg.txt",net0.n_4_7_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_3_zpos.txt",net0.n_4_7_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_3_zneg.txt",net0.n_4_7_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_4_local.txt",net0.n_4_7_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_4_xpos.txt",net0.n_4_7_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_4_xneg.txt",net0.n_4_7_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_4_ypos.txt",net0.n_4_7_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_4_yneg.txt",net0.n_4_7_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_4_zpos.txt",net0.n_4_7_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_4_zneg.txt",net0.n_4_7_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_4_xpos.txt",net0.n_4_7_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_4_xneg.txt",net0.n_4_7_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_4_ypos.txt",net0.n_4_7_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_4_yneg.txt",net0.n_4_7_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_4_zpos.txt",net0.n_4_7_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_4_zneg.txt",net0.n_4_7_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_4_xpos.txt",net0.n_4_7_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_4_xneg.txt",net0.n_4_7_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_4_ypos.txt",net0.n_4_7_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_4_yneg.txt",net0.n_4_7_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_4_zpos.txt",net0.n_4_7_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_4_zneg.txt",net0.n_4_7_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_5_local.txt",net0.n_4_7_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_5_xpos.txt",net0.n_4_7_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_5_xneg.txt",net0.n_4_7_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_5_ypos.txt",net0.n_4_7_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_5_yneg.txt",net0.n_4_7_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_5_zpos.txt",net0.n_4_7_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_5_zneg.txt",net0.n_4_7_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_5_xpos.txt",net0.n_4_7_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_5_xneg.txt",net0.n_4_7_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_5_ypos.txt",net0.n_4_7_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_5_yneg.txt",net0.n_4_7_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_5_zpos.txt",net0.n_4_7_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_5_zneg.txt",net0.n_4_7_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_5_xpos.txt",net0.n_4_7_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_5_xneg.txt",net0.n_4_7_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_5_ypos.txt",net0.n_4_7_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_5_yneg.txt",net0.n_4_7_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_5_zpos.txt",net0.n_4_7_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_5_zneg.txt",net0.n_4_7_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_6_local.txt",net0.n_4_7_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_6_xpos.txt",net0.n_4_7_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_6_xneg.txt",net0.n_4_7_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_6_ypos.txt",net0.n_4_7_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_6_yneg.txt",net0.n_4_7_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_6_zpos.txt",net0.n_4_7_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_6_zneg.txt",net0.n_4_7_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_6_xpos.txt",net0.n_4_7_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_6_xneg.txt",net0.n_4_7_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_6_ypos.txt",net0.n_4_7_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_6_yneg.txt",net0.n_4_7_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_6_zpos.txt",net0.n_4_7_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_6_zneg.txt",net0.n_4_7_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_6_xpos.txt",net0.n_4_7_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_6_xneg.txt",net0.n_4_7_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_6_ypos.txt",net0.n_4_7_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_6_yneg.txt",net0.n_4_7_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_6_zpos.txt",net0.n_4_7_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_6_zneg.txt",net0.n_4_7_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_7_local.txt",net0.n_4_7_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_7_xpos.txt",net0.n_4_7_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_7_xneg.txt",net0.n_4_7_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_7_ypos.txt",net0.n_4_7_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_7_yneg.txt",net0.n_4_7_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_7_zpos.txt",net0.n_4_7_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_4_7_7_zneg.txt",net0.n_4_7_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_7_xpos.txt",net0.n_4_7_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_7_xneg.txt",net0.n_4_7_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_7_ypos.txt",net0.n_4_7_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_7_yneg.txt",net0.n_4_7_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_7_zpos.txt",net0.n_4_7_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_4_7_7_zneg.txt",net0.n_4_7_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_7_xpos.txt",net0.n_4_7_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_7_xneg.txt",net0.n_4_7_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_7_ypos.txt",net0.n_4_7_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_7_yneg.txt",net0.n_4_7_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_7_zpos.txt",net0.n_4_7_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_4_7_7_zneg.txt",net0.n_4_7_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_0_local.txt",net0.n_5_0_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_0_xpos.txt",net0.n_5_0_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_0_xneg.txt",net0.n_5_0_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_0_ypos.txt",net0.n_5_0_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_0_yneg.txt",net0.n_5_0_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_0_zpos.txt",net0.n_5_0_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_0_zneg.txt",net0.n_5_0_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_0_xpos.txt",net0.n_5_0_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_0_xneg.txt",net0.n_5_0_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_0_ypos.txt",net0.n_5_0_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_0_yneg.txt",net0.n_5_0_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_0_zpos.txt",net0.n_5_0_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_0_zneg.txt",net0.n_5_0_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_0_xpos.txt",net0.n_5_0_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_0_xneg.txt",net0.n_5_0_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_0_ypos.txt",net0.n_5_0_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_0_yneg.txt",net0.n_5_0_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_0_zpos.txt",net0.n_5_0_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_0_zneg.txt",net0.n_5_0_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_1_local.txt",net0.n_5_0_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_1_xpos.txt",net0.n_5_0_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_1_xneg.txt",net0.n_5_0_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_1_ypos.txt",net0.n_5_0_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_1_yneg.txt",net0.n_5_0_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_1_zpos.txt",net0.n_5_0_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_1_zneg.txt",net0.n_5_0_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_1_xpos.txt",net0.n_5_0_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_1_xneg.txt",net0.n_5_0_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_1_ypos.txt",net0.n_5_0_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_1_yneg.txt",net0.n_5_0_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_1_zpos.txt",net0.n_5_0_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_1_zneg.txt",net0.n_5_0_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_1_xpos.txt",net0.n_5_0_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_1_xneg.txt",net0.n_5_0_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_1_ypos.txt",net0.n_5_0_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_1_yneg.txt",net0.n_5_0_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_1_zpos.txt",net0.n_5_0_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_1_zneg.txt",net0.n_5_0_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_2_local.txt",net0.n_5_0_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_2_xpos.txt",net0.n_5_0_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_2_xneg.txt",net0.n_5_0_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_2_ypos.txt",net0.n_5_0_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_2_yneg.txt",net0.n_5_0_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_2_zpos.txt",net0.n_5_0_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_2_zneg.txt",net0.n_5_0_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_2_xpos.txt",net0.n_5_0_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_2_xneg.txt",net0.n_5_0_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_2_ypos.txt",net0.n_5_0_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_2_yneg.txt",net0.n_5_0_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_2_zpos.txt",net0.n_5_0_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_2_zneg.txt",net0.n_5_0_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_2_xpos.txt",net0.n_5_0_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_2_xneg.txt",net0.n_5_0_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_2_ypos.txt",net0.n_5_0_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_2_yneg.txt",net0.n_5_0_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_2_zpos.txt",net0.n_5_0_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_2_zneg.txt",net0.n_5_0_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_3_local.txt",net0.n_5_0_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_3_xpos.txt",net0.n_5_0_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_3_xneg.txt",net0.n_5_0_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_3_ypos.txt",net0.n_5_0_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_3_yneg.txt",net0.n_5_0_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_3_zpos.txt",net0.n_5_0_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_3_zneg.txt",net0.n_5_0_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_3_xpos.txt",net0.n_5_0_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_3_xneg.txt",net0.n_5_0_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_3_ypos.txt",net0.n_5_0_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_3_yneg.txt",net0.n_5_0_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_3_zpos.txt",net0.n_5_0_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_3_zneg.txt",net0.n_5_0_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_3_xpos.txt",net0.n_5_0_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_3_xneg.txt",net0.n_5_0_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_3_ypos.txt",net0.n_5_0_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_3_yneg.txt",net0.n_5_0_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_3_zpos.txt",net0.n_5_0_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_3_zneg.txt",net0.n_5_0_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_4_local.txt",net0.n_5_0_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_4_xpos.txt",net0.n_5_0_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_4_xneg.txt",net0.n_5_0_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_4_ypos.txt",net0.n_5_0_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_4_yneg.txt",net0.n_5_0_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_4_zpos.txt",net0.n_5_0_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_4_zneg.txt",net0.n_5_0_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_4_xpos.txt",net0.n_5_0_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_4_xneg.txt",net0.n_5_0_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_4_ypos.txt",net0.n_5_0_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_4_yneg.txt",net0.n_5_0_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_4_zpos.txt",net0.n_5_0_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_4_zneg.txt",net0.n_5_0_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_4_xpos.txt",net0.n_5_0_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_4_xneg.txt",net0.n_5_0_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_4_ypos.txt",net0.n_5_0_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_4_yneg.txt",net0.n_5_0_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_4_zpos.txt",net0.n_5_0_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_4_zneg.txt",net0.n_5_0_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_5_local.txt",net0.n_5_0_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_5_xpos.txt",net0.n_5_0_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_5_xneg.txt",net0.n_5_0_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_5_ypos.txt",net0.n_5_0_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_5_yneg.txt",net0.n_5_0_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_5_zpos.txt",net0.n_5_0_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_5_zneg.txt",net0.n_5_0_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_5_xpos.txt",net0.n_5_0_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_5_xneg.txt",net0.n_5_0_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_5_ypos.txt",net0.n_5_0_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_5_yneg.txt",net0.n_5_0_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_5_zpos.txt",net0.n_5_0_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_5_zneg.txt",net0.n_5_0_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_5_xpos.txt",net0.n_5_0_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_5_xneg.txt",net0.n_5_0_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_5_ypos.txt",net0.n_5_0_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_5_yneg.txt",net0.n_5_0_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_5_zpos.txt",net0.n_5_0_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_5_zneg.txt",net0.n_5_0_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_6_local.txt",net0.n_5_0_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_6_xpos.txt",net0.n_5_0_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_6_xneg.txt",net0.n_5_0_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_6_ypos.txt",net0.n_5_0_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_6_yneg.txt",net0.n_5_0_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_6_zpos.txt",net0.n_5_0_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_6_zneg.txt",net0.n_5_0_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_6_xpos.txt",net0.n_5_0_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_6_xneg.txt",net0.n_5_0_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_6_ypos.txt",net0.n_5_0_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_6_yneg.txt",net0.n_5_0_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_6_zpos.txt",net0.n_5_0_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_6_zneg.txt",net0.n_5_0_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_6_xpos.txt",net0.n_5_0_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_6_xneg.txt",net0.n_5_0_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_6_ypos.txt",net0.n_5_0_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_6_yneg.txt",net0.n_5_0_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_6_zpos.txt",net0.n_5_0_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_6_zneg.txt",net0.n_5_0_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_7_local.txt",net0.n_5_0_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_7_xpos.txt",net0.n_5_0_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_7_xneg.txt",net0.n_5_0_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_7_ypos.txt",net0.n_5_0_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_7_yneg.txt",net0.n_5_0_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_7_zpos.txt",net0.n_5_0_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_0_7_zneg.txt",net0.n_5_0_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_7_xpos.txt",net0.n_5_0_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_7_xneg.txt",net0.n_5_0_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_7_ypos.txt",net0.n_5_0_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_7_yneg.txt",net0.n_5_0_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_7_zpos.txt",net0.n_5_0_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_0_7_zneg.txt",net0.n_5_0_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_7_xpos.txt",net0.n_5_0_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_7_xneg.txt",net0.n_5_0_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_7_ypos.txt",net0.n_5_0_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_7_yneg.txt",net0.n_5_0_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_7_zpos.txt",net0.n_5_0_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_0_7_zneg.txt",net0.n_5_0_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_0_local.txt",net0.n_5_1_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_0_xpos.txt",net0.n_5_1_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_0_xneg.txt",net0.n_5_1_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_0_ypos.txt",net0.n_5_1_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_0_yneg.txt",net0.n_5_1_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_0_zpos.txt",net0.n_5_1_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_0_zneg.txt",net0.n_5_1_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_0_xpos.txt",net0.n_5_1_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_0_xneg.txt",net0.n_5_1_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_0_ypos.txt",net0.n_5_1_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_0_yneg.txt",net0.n_5_1_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_0_zpos.txt",net0.n_5_1_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_0_zneg.txt",net0.n_5_1_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_0_xpos.txt",net0.n_5_1_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_0_xneg.txt",net0.n_5_1_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_0_ypos.txt",net0.n_5_1_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_0_yneg.txt",net0.n_5_1_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_0_zpos.txt",net0.n_5_1_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_0_zneg.txt",net0.n_5_1_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_1_local.txt",net0.n_5_1_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_1_xpos.txt",net0.n_5_1_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_1_xneg.txt",net0.n_5_1_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_1_ypos.txt",net0.n_5_1_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_1_yneg.txt",net0.n_5_1_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_1_zpos.txt",net0.n_5_1_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_1_zneg.txt",net0.n_5_1_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_1_xpos.txt",net0.n_5_1_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_1_xneg.txt",net0.n_5_1_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_1_ypos.txt",net0.n_5_1_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_1_yneg.txt",net0.n_5_1_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_1_zpos.txt",net0.n_5_1_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_1_zneg.txt",net0.n_5_1_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_1_xpos.txt",net0.n_5_1_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_1_xneg.txt",net0.n_5_1_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_1_ypos.txt",net0.n_5_1_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_1_yneg.txt",net0.n_5_1_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_1_zpos.txt",net0.n_5_1_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_1_zneg.txt",net0.n_5_1_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_2_local.txt",net0.n_5_1_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_2_xpos.txt",net0.n_5_1_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_2_xneg.txt",net0.n_5_1_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_2_ypos.txt",net0.n_5_1_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_2_yneg.txt",net0.n_5_1_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_2_zpos.txt",net0.n_5_1_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_2_zneg.txt",net0.n_5_1_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_2_xpos.txt",net0.n_5_1_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_2_xneg.txt",net0.n_5_1_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_2_ypos.txt",net0.n_5_1_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_2_yneg.txt",net0.n_5_1_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_2_zpos.txt",net0.n_5_1_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_2_zneg.txt",net0.n_5_1_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_2_xpos.txt",net0.n_5_1_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_2_xneg.txt",net0.n_5_1_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_2_ypos.txt",net0.n_5_1_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_2_yneg.txt",net0.n_5_1_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_2_zpos.txt",net0.n_5_1_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_2_zneg.txt",net0.n_5_1_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_3_local.txt",net0.n_5_1_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_3_xpos.txt",net0.n_5_1_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_3_xneg.txt",net0.n_5_1_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_3_ypos.txt",net0.n_5_1_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_3_yneg.txt",net0.n_5_1_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_3_zpos.txt",net0.n_5_1_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_3_zneg.txt",net0.n_5_1_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_3_xpos.txt",net0.n_5_1_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_3_xneg.txt",net0.n_5_1_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_3_ypos.txt",net0.n_5_1_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_3_yneg.txt",net0.n_5_1_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_3_zpos.txt",net0.n_5_1_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_3_zneg.txt",net0.n_5_1_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_3_xpos.txt",net0.n_5_1_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_3_xneg.txt",net0.n_5_1_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_3_ypos.txt",net0.n_5_1_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_3_yneg.txt",net0.n_5_1_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_3_zpos.txt",net0.n_5_1_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_3_zneg.txt",net0.n_5_1_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_4_local.txt",net0.n_5_1_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_4_xpos.txt",net0.n_5_1_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_4_xneg.txt",net0.n_5_1_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_4_ypos.txt",net0.n_5_1_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_4_yneg.txt",net0.n_5_1_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_4_zpos.txt",net0.n_5_1_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_4_zneg.txt",net0.n_5_1_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_4_xpos.txt",net0.n_5_1_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_4_xneg.txt",net0.n_5_1_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_4_ypos.txt",net0.n_5_1_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_4_yneg.txt",net0.n_5_1_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_4_zpos.txt",net0.n_5_1_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_4_zneg.txt",net0.n_5_1_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_4_xpos.txt",net0.n_5_1_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_4_xneg.txt",net0.n_5_1_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_4_ypos.txt",net0.n_5_1_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_4_yneg.txt",net0.n_5_1_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_4_zpos.txt",net0.n_5_1_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_4_zneg.txt",net0.n_5_1_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_5_local.txt",net0.n_5_1_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_5_xpos.txt",net0.n_5_1_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_5_xneg.txt",net0.n_5_1_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_5_ypos.txt",net0.n_5_1_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_5_yneg.txt",net0.n_5_1_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_5_zpos.txt",net0.n_5_1_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_5_zneg.txt",net0.n_5_1_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_5_xpos.txt",net0.n_5_1_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_5_xneg.txt",net0.n_5_1_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_5_ypos.txt",net0.n_5_1_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_5_yneg.txt",net0.n_5_1_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_5_zpos.txt",net0.n_5_1_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_5_zneg.txt",net0.n_5_1_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_5_xpos.txt",net0.n_5_1_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_5_xneg.txt",net0.n_5_1_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_5_ypos.txt",net0.n_5_1_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_5_yneg.txt",net0.n_5_1_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_5_zpos.txt",net0.n_5_1_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_5_zneg.txt",net0.n_5_1_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_6_local.txt",net0.n_5_1_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_6_xpos.txt",net0.n_5_1_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_6_xneg.txt",net0.n_5_1_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_6_ypos.txt",net0.n_5_1_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_6_yneg.txt",net0.n_5_1_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_6_zpos.txt",net0.n_5_1_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_6_zneg.txt",net0.n_5_1_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_6_xpos.txt",net0.n_5_1_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_6_xneg.txt",net0.n_5_1_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_6_ypos.txt",net0.n_5_1_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_6_yneg.txt",net0.n_5_1_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_6_zpos.txt",net0.n_5_1_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_6_zneg.txt",net0.n_5_1_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_6_xpos.txt",net0.n_5_1_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_6_xneg.txt",net0.n_5_1_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_6_ypos.txt",net0.n_5_1_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_6_yneg.txt",net0.n_5_1_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_6_zpos.txt",net0.n_5_1_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_6_zneg.txt",net0.n_5_1_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_7_local.txt",net0.n_5_1_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_7_xpos.txt",net0.n_5_1_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_7_xneg.txt",net0.n_5_1_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_7_ypos.txt",net0.n_5_1_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_7_yneg.txt",net0.n_5_1_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_7_zpos.txt",net0.n_5_1_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_1_7_zneg.txt",net0.n_5_1_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_7_xpos.txt",net0.n_5_1_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_7_xneg.txt",net0.n_5_1_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_7_ypos.txt",net0.n_5_1_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_7_yneg.txt",net0.n_5_1_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_7_zpos.txt",net0.n_5_1_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_1_7_zneg.txt",net0.n_5_1_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_7_xpos.txt",net0.n_5_1_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_7_xneg.txt",net0.n_5_1_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_7_ypos.txt",net0.n_5_1_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_7_yneg.txt",net0.n_5_1_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_7_zpos.txt",net0.n_5_1_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_1_7_zneg.txt",net0.n_5_1_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_0_local.txt",net0.n_5_2_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_0_xpos.txt",net0.n_5_2_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_0_xneg.txt",net0.n_5_2_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_0_ypos.txt",net0.n_5_2_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_0_yneg.txt",net0.n_5_2_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_0_zpos.txt",net0.n_5_2_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_0_zneg.txt",net0.n_5_2_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_0_xpos.txt",net0.n_5_2_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_0_xneg.txt",net0.n_5_2_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_0_ypos.txt",net0.n_5_2_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_0_yneg.txt",net0.n_5_2_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_0_zpos.txt",net0.n_5_2_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_0_zneg.txt",net0.n_5_2_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_0_xpos.txt",net0.n_5_2_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_0_xneg.txt",net0.n_5_2_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_0_ypos.txt",net0.n_5_2_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_0_yneg.txt",net0.n_5_2_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_0_zpos.txt",net0.n_5_2_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_0_zneg.txt",net0.n_5_2_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_1_local.txt",net0.n_5_2_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_1_xpos.txt",net0.n_5_2_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_1_xneg.txt",net0.n_5_2_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_1_ypos.txt",net0.n_5_2_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_1_yneg.txt",net0.n_5_2_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_1_zpos.txt",net0.n_5_2_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_1_zneg.txt",net0.n_5_2_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_1_xpos.txt",net0.n_5_2_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_1_xneg.txt",net0.n_5_2_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_1_ypos.txt",net0.n_5_2_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_1_yneg.txt",net0.n_5_2_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_1_zpos.txt",net0.n_5_2_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_1_zneg.txt",net0.n_5_2_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_1_xpos.txt",net0.n_5_2_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_1_xneg.txt",net0.n_5_2_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_1_ypos.txt",net0.n_5_2_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_1_yneg.txt",net0.n_5_2_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_1_zpos.txt",net0.n_5_2_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_1_zneg.txt",net0.n_5_2_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_2_local.txt",net0.n_5_2_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_2_xpos.txt",net0.n_5_2_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_2_xneg.txt",net0.n_5_2_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_2_ypos.txt",net0.n_5_2_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_2_yneg.txt",net0.n_5_2_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_2_zpos.txt",net0.n_5_2_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_2_zneg.txt",net0.n_5_2_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_2_xpos.txt",net0.n_5_2_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_2_xneg.txt",net0.n_5_2_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_2_ypos.txt",net0.n_5_2_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_2_yneg.txt",net0.n_5_2_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_2_zpos.txt",net0.n_5_2_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_2_zneg.txt",net0.n_5_2_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_2_xpos.txt",net0.n_5_2_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_2_xneg.txt",net0.n_5_2_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_2_ypos.txt",net0.n_5_2_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_2_yneg.txt",net0.n_5_2_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_2_zpos.txt",net0.n_5_2_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_2_zneg.txt",net0.n_5_2_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_3_local.txt",net0.n_5_2_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_3_xpos.txt",net0.n_5_2_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_3_xneg.txt",net0.n_5_2_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_3_ypos.txt",net0.n_5_2_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_3_yneg.txt",net0.n_5_2_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_3_zpos.txt",net0.n_5_2_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_3_zneg.txt",net0.n_5_2_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_3_xpos.txt",net0.n_5_2_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_3_xneg.txt",net0.n_5_2_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_3_ypos.txt",net0.n_5_2_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_3_yneg.txt",net0.n_5_2_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_3_zpos.txt",net0.n_5_2_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_3_zneg.txt",net0.n_5_2_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_3_xpos.txt",net0.n_5_2_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_3_xneg.txt",net0.n_5_2_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_3_ypos.txt",net0.n_5_2_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_3_yneg.txt",net0.n_5_2_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_3_zpos.txt",net0.n_5_2_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_3_zneg.txt",net0.n_5_2_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_4_local.txt",net0.n_5_2_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_4_xpos.txt",net0.n_5_2_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_4_xneg.txt",net0.n_5_2_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_4_ypos.txt",net0.n_5_2_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_4_yneg.txt",net0.n_5_2_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_4_zpos.txt",net0.n_5_2_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_4_zneg.txt",net0.n_5_2_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_4_xpos.txt",net0.n_5_2_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_4_xneg.txt",net0.n_5_2_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_4_ypos.txt",net0.n_5_2_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_4_yneg.txt",net0.n_5_2_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_4_zpos.txt",net0.n_5_2_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_4_zneg.txt",net0.n_5_2_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_4_xpos.txt",net0.n_5_2_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_4_xneg.txt",net0.n_5_2_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_4_ypos.txt",net0.n_5_2_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_4_yneg.txt",net0.n_5_2_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_4_zpos.txt",net0.n_5_2_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_4_zneg.txt",net0.n_5_2_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_5_local.txt",net0.n_5_2_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_5_xpos.txt",net0.n_5_2_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_5_xneg.txt",net0.n_5_2_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_5_ypos.txt",net0.n_5_2_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_5_yneg.txt",net0.n_5_2_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_5_zpos.txt",net0.n_5_2_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_5_zneg.txt",net0.n_5_2_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_5_xpos.txt",net0.n_5_2_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_5_xneg.txt",net0.n_5_2_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_5_ypos.txt",net0.n_5_2_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_5_yneg.txt",net0.n_5_2_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_5_zpos.txt",net0.n_5_2_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_5_zneg.txt",net0.n_5_2_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_5_xpos.txt",net0.n_5_2_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_5_xneg.txt",net0.n_5_2_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_5_ypos.txt",net0.n_5_2_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_5_yneg.txt",net0.n_5_2_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_5_zpos.txt",net0.n_5_2_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_5_zneg.txt",net0.n_5_2_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_6_local.txt",net0.n_5_2_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_6_xpos.txt",net0.n_5_2_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_6_xneg.txt",net0.n_5_2_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_6_ypos.txt",net0.n_5_2_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_6_yneg.txt",net0.n_5_2_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_6_zpos.txt",net0.n_5_2_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_6_zneg.txt",net0.n_5_2_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_6_xpos.txt",net0.n_5_2_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_6_xneg.txt",net0.n_5_2_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_6_ypos.txt",net0.n_5_2_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_6_yneg.txt",net0.n_5_2_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_6_zpos.txt",net0.n_5_2_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_6_zneg.txt",net0.n_5_2_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_6_xpos.txt",net0.n_5_2_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_6_xneg.txt",net0.n_5_2_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_6_ypos.txt",net0.n_5_2_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_6_yneg.txt",net0.n_5_2_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_6_zpos.txt",net0.n_5_2_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_6_zneg.txt",net0.n_5_2_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_7_local.txt",net0.n_5_2_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_7_xpos.txt",net0.n_5_2_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_7_xneg.txt",net0.n_5_2_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_7_ypos.txt",net0.n_5_2_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_7_yneg.txt",net0.n_5_2_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_7_zpos.txt",net0.n_5_2_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_2_7_zneg.txt",net0.n_5_2_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_7_xpos.txt",net0.n_5_2_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_7_xneg.txt",net0.n_5_2_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_7_ypos.txt",net0.n_5_2_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_7_yneg.txt",net0.n_5_2_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_7_zpos.txt",net0.n_5_2_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_2_7_zneg.txt",net0.n_5_2_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_7_xpos.txt",net0.n_5_2_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_7_xneg.txt",net0.n_5_2_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_7_ypos.txt",net0.n_5_2_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_7_yneg.txt",net0.n_5_2_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_7_zpos.txt",net0.n_5_2_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_2_7_zneg.txt",net0.n_5_2_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_0_local.txt",net0.n_5_3_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_0_xpos.txt",net0.n_5_3_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_0_xneg.txt",net0.n_5_3_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_0_ypos.txt",net0.n_5_3_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_0_yneg.txt",net0.n_5_3_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_0_zpos.txt",net0.n_5_3_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_0_zneg.txt",net0.n_5_3_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_0_xpos.txt",net0.n_5_3_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_0_xneg.txt",net0.n_5_3_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_0_ypos.txt",net0.n_5_3_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_0_yneg.txt",net0.n_5_3_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_0_zpos.txt",net0.n_5_3_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_0_zneg.txt",net0.n_5_3_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_0_xpos.txt",net0.n_5_3_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_0_xneg.txt",net0.n_5_3_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_0_ypos.txt",net0.n_5_3_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_0_yneg.txt",net0.n_5_3_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_0_zpos.txt",net0.n_5_3_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_0_zneg.txt",net0.n_5_3_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_1_local.txt",net0.n_5_3_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_1_xpos.txt",net0.n_5_3_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_1_xneg.txt",net0.n_5_3_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_1_ypos.txt",net0.n_5_3_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_1_yneg.txt",net0.n_5_3_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_1_zpos.txt",net0.n_5_3_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_1_zneg.txt",net0.n_5_3_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_1_xpos.txt",net0.n_5_3_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_1_xneg.txt",net0.n_5_3_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_1_ypos.txt",net0.n_5_3_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_1_yneg.txt",net0.n_5_3_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_1_zpos.txt",net0.n_5_3_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_1_zneg.txt",net0.n_5_3_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_1_xpos.txt",net0.n_5_3_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_1_xneg.txt",net0.n_5_3_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_1_ypos.txt",net0.n_5_3_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_1_yneg.txt",net0.n_5_3_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_1_zpos.txt",net0.n_5_3_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_1_zneg.txt",net0.n_5_3_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_2_local.txt",net0.n_5_3_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_2_xpos.txt",net0.n_5_3_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_2_xneg.txt",net0.n_5_3_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_2_ypos.txt",net0.n_5_3_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_2_yneg.txt",net0.n_5_3_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_2_zpos.txt",net0.n_5_3_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_2_zneg.txt",net0.n_5_3_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_2_xpos.txt",net0.n_5_3_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_2_xneg.txt",net0.n_5_3_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_2_ypos.txt",net0.n_5_3_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_2_yneg.txt",net0.n_5_3_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_2_zpos.txt",net0.n_5_3_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_2_zneg.txt",net0.n_5_3_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_2_xpos.txt",net0.n_5_3_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_2_xneg.txt",net0.n_5_3_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_2_ypos.txt",net0.n_5_3_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_2_yneg.txt",net0.n_5_3_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_2_zpos.txt",net0.n_5_3_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_2_zneg.txt",net0.n_5_3_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_3_local.txt",net0.n_5_3_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_3_xpos.txt",net0.n_5_3_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_3_xneg.txt",net0.n_5_3_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_3_ypos.txt",net0.n_5_3_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_3_yneg.txt",net0.n_5_3_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_3_zpos.txt",net0.n_5_3_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_3_zneg.txt",net0.n_5_3_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_3_xpos.txt",net0.n_5_3_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_3_xneg.txt",net0.n_5_3_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_3_ypos.txt",net0.n_5_3_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_3_yneg.txt",net0.n_5_3_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_3_zpos.txt",net0.n_5_3_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_3_zneg.txt",net0.n_5_3_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_3_xpos.txt",net0.n_5_3_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_3_xneg.txt",net0.n_5_3_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_3_ypos.txt",net0.n_5_3_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_3_yneg.txt",net0.n_5_3_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_3_zpos.txt",net0.n_5_3_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_3_zneg.txt",net0.n_5_3_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_4_local.txt",net0.n_5_3_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_4_xpos.txt",net0.n_5_3_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_4_xneg.txt",net0.n_5_3_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_4_ypos.txt",net0.n_5_3_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_4_yneg.txt",net0.n_5_3_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_4_zpos.txt",net0.n_5_3_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_4_zneg.txt",net0.n_5_3_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_4_xpos.txt",net0.n_5_3_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_4_xneg.txt",net0.n_5_3_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_4_ypos.txt",net0.n_5_3_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_4_yneg.txt",net0.n_5_3_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_4_zpos.txt",net0.n_5_3_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_4_zneg.txt",net0.n_5_3_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_4_xpos.txt",net0.n_5_3_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_4_xneg.txt",net0.n_5_3_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_4_ypos.txt",net0.n_5_3_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_4_yneg.txt",net0.n_5_3_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_4_zpos.txt",net0.n_5_3_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_4_zneg.txt",net0.n_5_3_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_5_local.txt",net0.n_5_3_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_5_xpos.txt",net0.n_5_3_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_5_xneg.txt",net0.n_5_3_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_5_ypos.txt",net0.n_5_3_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_5_yneg.txt",net0.n_5_3_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_5_zpos.txt",net0.n_5_3_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_5_zneg.txt",net0.n_5_3_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_5_xpos.txt",net0.n_5_3_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_5_xneg.txt",net0.n_5_3_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_5_ypos.txt",net0.n_5_3_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_5_yneg.txt",net0.n_5_3_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_5_zpos.txt",net0.n_5_3_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_5_zneg.txt",net0.n_5_3_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_5_xpos.txt",net0.n_5_3_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_5_xneg.txt",net0.n_5_3_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_5_ypos.txt",net0.n_5_3_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_5_yneg.txt",net0.n_5_3_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_5_zpos.txt",net0.n_5_3_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_5_zneg.txt",net0.n_5_3_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_6_local.txt",net0.n_5_3_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_6_xpos.txt",net0.n_5_3_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_6_xneg.txt",net0.n_5_3_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_6_ypos.txt",net0.n_5_3_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_6_yneg.txt",net0.n_5_3_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_6_zpos.txt",net0.n_5_3_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_6_zneg.txt",net0.n_5_3_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_6_xpos.txt",net0.n_5_3_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_6_xneg.txt",net0.n_5_3_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_6_ypos.txt",net0.n_5_3_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_6_yneg.txt",net0.n_5_3_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_6_zpos.txt",net0.n_5_3_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_6_zneg.txt",net0.n_5_3_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_6_xpos.txt",net0.n_5_3_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_6_xneg.txt",net0.n_5_3_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_6_ypos.txt",net0.n_5_3_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_6_yneg.txt",net0.n_5_3_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_6_zpos.txt",net0.n_5_3_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_6_zneg.txt",net0.n_5_3_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_7_local.txt",net0.n_5_3_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_7_xpos.txt",net0.n_5_3_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_7_xneg.txt",net0.n_5_3_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_7_ypos.txt",net0.n_5_3_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_7_yneg.txt",net0.n_5_3_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_7_zpos.txt",net0.n_5_3_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_3_7_zneg.txt",net0.n_5_3_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_7_xpos.txt",net0.n_5_3_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_7_xneg.txt",net0.n_5_3_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_7_ypos.txt",net0.n_5_3_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_7_yneg.txt",net0.n_5_3_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_7_zpos.txt",net0.n_5_3_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_3_7_zneg.txt",net0.n_5_3_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_7_xpos.txt",net0.n_5_3_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_7_xneg.txt",net0.n_5_3_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_7_ypos.txt",net0.n_5_3_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_7_yneg.txt",net0.n_5_3_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_7_zpos.txt",net0.n_5_3_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_3_7_zneg.txt",net0.n_5_3_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_0_local.txt",net0.n_5_4_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_0_xpos.txt",net0.n_5_4_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_0_xneg.txt",net0.n_5_4_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_0_ypos.txt",net0.n_5_4_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_0_yneg.txt",net0.n_5_4_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_0_zpos.txt",net0.n_5_4_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_0_zneg.txt",net0.n_5_4_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_0_xpos.txt",net0.n_5_4_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_0_xneg.txt",net0.n_5_4_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_0_ypos.txt",net0.n_5_4_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_0_yneg.txt",net0.n_5_4_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_0_zpos.txt",net0.n_5_4_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_0_zneg.txt",net0.n_5_4_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_0_xpos.txt",net0.n_5_4_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_0_xneg.txt",net0.n_5_4_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_0_ypos.txt",net0.n_5_4_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_0_yneg.txt",net0.n_5_4_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_0_zpos.txt",net0.n_5_4_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_0_zneg.txt",net0.n_5_4_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_1_local.txt",net0.n_5_4_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_1_xpos.txt",net0.n_5_4_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_1_xneg.txt",net0.n_5_4_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_1_ypos.txt",net0.n_5_4_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_1_yneg.txt",net0.n_5_4_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_1_zpos.txt",net0.n_5_4_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_1_zneg.txt",net0.n_5_4_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_1_xpos.txt",net0.n_5_4_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_1_xneg.txt",net0.n_5_4_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_1_ypos.txt",net0.n_5_4_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_1_yneg.txt",net0.n_5_4_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_1_zpos.txt",net0.n_5_4_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_1_zneg.txt",net0.n_5_4_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_1_xpos.txt",net0.n_5_4_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_1_xneg.txt",net0.n_5_4_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_1_ypos.txt",net0.n_5_4_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_1_yneg.txt",net0.n_5_4_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_1_zpos.txt",net0.n_5_4_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_1_zneg.txt",net0.n_5_4_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_2_local.txt",net0.n_5_4_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_2_xpos.txt",net0.n_5_4_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_2_xneg.txt",net0.n_5_4_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_2_ypos.txt",net0.n_5_4_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_2_yneg.txt",net0.n_5_4_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_2_zpos.txt",net0.n_5_4_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_2_zneg.txt",net0.n_5_4_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_2_xpos.txt",net0.n_5_4_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_2_xneg.txt",net0.n_5_4_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_2_ypos.txt",net0.n_5_4_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_2_yneg.txt",net0.n_5_4_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_2_zpos.txt",net0.n_5_4_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_2_zneg.txt",net0.n_5_4_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_2_xpos.txt",net0.n_5_4_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_2_xneg.txt",net0.n_5_4_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_2_ypos.txt",net0.n_5_4_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_2_yneg.txt",net0.n_5_4_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_2_zpos.txt",net0.n_5_4_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_2_zneg.txt",net0.n_5_4_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_3_local.txt",net0.n_5_4_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_3_xpos.txt",net0.n_5_4_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_3_xneg.txt",net0.n_5_4_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_3_ypos.txt",net0.n_5_4_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_3_yneg.txt",net0.n_5_4_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_3_zpos.txt",net0.n_5_4_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_3_zneg.txt",net0.n_5_4_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_3_xpos.txt",net0.n_5_4_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_3_xneg.txt",net0.n_5_4_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_3_ypos.txt",net0.n_5_4_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_3_yneg.txt",net0.n_5_4_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_3_zpos.txt",net0.n_5_4_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_3_zneg.txt",net0.n_5_4_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_3_xpos.txt",net0.n_5_4_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_3_xneg.txt",net0.n_5_4_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_3_ypos.txt",net0.n_5_4_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_3_yneg.txt",net0.n_5_4_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_3_zpos.txt",net0.n_5_4_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_3_zneg.txt",net0.n_5_4_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_4_local.txt",net0.n_5_4_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_4_xpos.txt",net0.n_5_4_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_4_xneg.txt",net0.n_5_4_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_4_ypos.txt",net0.n_5_4_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_4_yneg.txt",net0.n_5_4_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_4_zpos.txt",net0.n_5_4_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_4_zneg.txt",net0.n_5_4_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_4_xpos.txt",net0.n_5_4_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_4_xneg.txt",net0.n_5_4_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_4_ypos.txt",net0.n_5_4_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_4_yneg.txt",net0.n_5_4_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_4_zpos.txt",net0.n_5_4_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_4_zneg.txt",net0.n_5_4_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_4_xpos.txt",net0.n_5_4_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_4_xneg.txt",net0.n_5_4_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_4_ypos.txt",net0.n_5_4_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_4_yneg.txt",net0.n_5_4_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_4_zpos.txt",net0.n_5_4_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_4_zneg.txt",net0.n_5_4_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_5_local.txt",net0.n_5_4_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_5_xpos.txt",net0.n_5_4_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_5_xneg.txt",net0.n_5_4_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_5_ypos.txt",net0.n_5_4_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_5_yneg.txt",net0.n_5_4_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_5_zpos.txt",net0.n_5_4_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_5_zneg.txt",net0.n_5_4_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_5_xpos.txt",net0.n_5_4_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_5_xneg.txt",net0.n_5_4_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_5_ypos.txt",net0.n_5_4_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_5_yneg.txt",net0.n_5_4_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_5_zpos.txt",net0.n_5_4_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_5_zneg.txt",net0.n_5_4_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_5_xpos.txt",net0.n_5_4_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_5_xneg.txt",net0.n_5_4_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_5_ypos.txt",net0.n_5_4_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_5_yneg.txt",net0.n_5_4_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_5_zpos.txt",net0.n_5_4_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_5_zneg.txt",net0.n_5_4_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_6_local.txt",net0.n_5_4_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_6_xpos.txt",net0.n_5_4_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_6_xneg.txt",net0.n_5_4_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_6_ypos.txt",net0.n_5_4_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_6_yneg.txt",net0.n_5_4_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_6_zpos.txt",net0.n_5_4_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_6_zneg.txt",net0.n_5_4_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_6_xpos.txt",net0.n_5_4_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_6_xneg.txt",net0.n_5_4_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_6_ypos.txt",net0.n_5_4_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_6_yneg.txt",net0.n_5_4_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_6_zpos.txt",net0.n_5_4_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_6_zneg.txt",net0.n_5_4_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_6_xpos.txt",net0.n_5_4_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_6_xneg.txt",net0.n_5_4_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_6_ypos.txt",net0.n_5_4_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_6_yneg.txt",net0.n_5_4_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_6_zpos.txt",net0.n_5_4_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_6_zneg.txt",net0.n_5_4_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_7_local.txt",net0.n_5_4_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_7_xpos.txt",net0.n_5_4_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_7_xneg.txt",net0.n_5_4_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_7_ypos.txt",net0.n_5_4_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_7_yneg.txt",net0.n_5_4_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_7_zpos.txt",net0.n_5_4_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_4_7_zneg.txt",net0.n_5_4_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_7_xpos.txt",net0.n_5_4_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_7_xneg.txt",net0.n_5_4_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_7_ypos.txt",net0.n_5_4_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_7_yneg.txt",net0.n_5_4_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_7_zpos.txt",net0.n_5_4_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_4_7_zneg.txt",net0.n_5_4_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_7_xpos.txt",net0.n_5_4_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_7_xneg.txt",net0.n_5_4_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_7_ypos.txt",net0.n_5_4_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_7_yneg.txt",net0.n_5_4_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_7_zpos.txt",net0.n_5_4_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_4_7_zneg.txt",net0.n_5_4_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_0_local.txt",net0.n_5_5_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_0_xpos.txt",net0.n_5_5_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_0_xneg.txt",net0.n_5_5_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_0_ypos.txt",net0.n_5_5_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_0_yneg.txt",net0.n_5_5_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_0_zpos.txt",net0.n_5_5_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_0_zneg.txt",net0.n_5_5_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_0_xpos.txt",net0.n_5_5_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_0_xneg.txt",net0.n_5_5_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_0_ypos.txt",net0.n_5_5_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_0_yneg.txt",net0.n_5_5_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_0_zpos.txt",net0.n_5_5_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_0_zneg.txt",net0.n_5_5_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_0_xpos.txt",net0.n_5_5_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_0_xneg.txt",net0.n_5_5_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_0_ypos.txt",net0.n_5_5_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_0_yneg.txt",net0.n_5_5_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_0_zpos.txt",net0.n_5_5_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_0_zneg.txt",net0.n_5_5_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_1_local.txt",net0.n_5_5_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_1_xpos.txt",net0.n_5_5_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_1_xneg.txt",net0.n_5_5_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_1_ypos.txt",net0.n_5_5_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_1_yneg.txt",net0.n_5_5_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_1_zpos.txt",net0.n_5_5_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_1_zneg.txt",net0.n_5_5_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_1_xpos.txt",net0.n_5_5_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_1_xneg.txt",net0.n_5_5_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_1_ypos.txt",net0.n_5_5_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_1_yneg.txt",net0.n_5_5_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_1_zpos.txt",net0.n_5_5_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_1_zneg.txt",net0.n_5_5_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_1_xpos.txt",net0.n_5_5_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_1_xneg.txt",net0.n_5_5_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_1_ypos.txt",net0.n_5_5_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_1_yneg.txt",net0.n_5_5_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_1_zpos.txt",net0.n_5_5_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_1_zneg.txt",net0.n_5_5_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_2_local.txt",net0.n_5_5_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_2_xpos.txt",net0.n_5_5_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_2_xneg.txt",net0.n_5_5_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_2_ypos.txt",net0.n_5_5_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_2_yneg.txt",net0.n_5_5_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_2_zpos.txt",net0.n_5_5_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_2_zneg.txt",net0.n_5_5_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_2_xpos.txt",net0.n_5_5_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_2_xneg.txt",net0.n_5_5_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_2_ypos.txt",net0.n_5_5_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_2_yneg.txt",net0.n_5_5_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_2_zpos.txt",net0.n_5_5_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_2_zneg.txt",net0.n_5_5_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_2_xpos.txt",net0.n_5_5_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_2_xneg.txt",net0.n_5_5_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_2_ypos.txt",net0.n_5_5_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_2_yneg.txt",net0.n_5_5_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_2_zpos.txt",net0.n_5_5_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_2_zneg.txt",net0.n_5_5_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_3_local.txt",net0.n_5_5_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_3_xpos.txt",net0.n_5_5_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_3_xneg.txt",net0.n_5_5_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_3_ypos.txt",net0.n_5_5_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_3_yneg.txt",net0.n_5_5_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_3_zpos.txt",net0.n_5_5_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_3_zneg.txt",net0.n_5_5_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_3_xpos.txt",net0.n_5_5_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_3_xneg.txt",net0.n_5_5_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_3_ypos.txt",net0.n_5_5_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_3_yneg.txt",net0.n_5_5_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_3_zpos.txt",net0.n_5_5_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_3_zneg.txt",net0.n_5_5_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_3_xpos.txt",net0.n_5_5_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_3_xneg.txt",net0.n_5_5_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_3_ypos.txt",net0.n_5_5_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_3_yneg.txt",net0.n_5_5_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_3_zpos.txt",net0.n_5_5_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_3_zneg.txt",net0.n_5_5_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_4_local.txt",net0.n_5_5_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_4_xpos.txt",net0.n_5_5_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_4_xneg.txt",net0.n_5_5_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_4_ypos.txt",net0.n_5_5_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_4_yneg.txt",net0.n_5_5_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_4_zpos.txt",net0.n_5_5_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_4_zneg.txt",net0.n_5_5_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_4_xpos.txt",net0.n_5_5_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_4_xneg.txt",net0.n_5_5_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_4_ypos.txt",net0.n_5_5_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_4_yneg.txt",net0.n_5_5_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_4_zpos.txt",net0.n_5_5_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_4_zneg.txt",net0.n_5_5_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_4_xpos.txt",net0.n_5_5_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_4_xneg.txt",net0.n_5_5_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_4_ypos.txt",net0.n_5_5_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_4_yneg.txt",net0.n_5_5_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_4_zpos.txt",net0.n_5_5_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_4_zneg.txt",net0.n_5_5_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_5_local.txt",net0.n_5_5_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_5_xpos.txt",net0.n_5_5_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_5_xneg.txt",net0.n_5_5_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_5_ypos.txt",net0.n_5_5_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_5_yneg.txt",net0.n_5_5_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_5_zpos.txt",net0.n_5_5_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_5_zneg.txt",net0.n_5_5_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_5_xpos.txt",net0.n_5_5_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_5_xneg.txt",net0.n_5_5_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_5_ypos.txt",net0.n_5_5_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_5_yneg.txt",net0.n_5_5_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_5_zpos.txt",net0.n_5_5_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_5_zneg.txt",net0.n_5_5_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_5_xpos.txt",net0.n_5_5_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_5_xneg.txt",net0.n_5_5_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_5_ypos.txt",net0.n_5_5_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_5_yneg.txt",net0.n_5_5_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_5_zpos.txt",net0.n_5_5_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_5_zneg.txt",net0.n_5_5_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_6_local.txt",net0.n_5_5_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_6_xpos.txt",net0.n_5_5_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_6_xneg.txt",net0.n_5_5_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_6_ypos.txt",net0.n_5_5_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_6_yneg.txt",net0.n_5_5_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_6_zpos.txt",net0.n_5_5_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_6_zneg.txt",net0.n_5_5_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_6_xpos.txt",net0.n_5_5_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_6_xneg.txt",net0.n_5_5_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_6_ypos.txt",net0.n_5_5_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_6_yneg.txt",net0.n_5_5_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_6_zpos.txt",net0.n_5_5_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_6_zneg.txt",net0.n_5_5_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_6_xpos.txt",net0.n_5_5_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_6_xneg.txt",net0.n_5_5_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_6_ypos.txt",net0.n_5_5_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_6_yneg.txt",net0.n_5_5_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_6_zpos.txt",net0.n_5_5_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_6_zneg.txt",net0.n_5_5_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_7_local.txt",net0.n_5_5_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_7_xpos.txt",net0.n_5_5_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_7_xneg.txt",net0.n_5_5_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_7_ypos.txt",net0.n_5_5_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_7_yneg.txt",net0.n_5_5_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_7_zpos.txt",net0.n_5_5_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_5_7_zneg.txt",net0.n_5_5_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_7_xpos.txt",net0.n_5_5_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_7_xneg.txt",net0.n_5_5_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_7_ypos.txt",net0.n_5_5_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_7_yneg.txt",net0.n_5_5_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_7_zpos.txt",net0.n_5_5_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_5_7_zneg.txt",net0.n_5_5_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_7_xpos.txt",net0.n_5_5_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_7_xneg.txt",net0.n_5_5_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_7_ypos.txt",net0.n_5_5_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_7_yneg.txt",net0.n_5_5_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_7_zpos.txt",net0.n_5_5_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_5_7_zneg.txt",net0.n_5_5_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_0_local.txt",net0.n_5_6_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_0_xpos.txt",net0.n_5_6_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_0_xneg.txt",net0.n_5_6_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_0_ypos.txt",net0.n_5_6_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_0_yneg.txt",net0.n_5_6_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_0_zpos.txt",net0.n_5_6_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_0_zneg.txt",net0.n_5_6_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_0_xpos.txt",net0.n_5_6_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_0_xneg.txt",net0.n_5_6_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_0_ypos.txt",net0.n_5_6_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_0_yneg.txt",net0.n_5_6_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_0_zpos.txt",net0.n_5_6_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_0_zneg.txt",net0.n_5_6_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_0_xpos.txt",net0.n_5_6_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_0_xneg.txt",net0.n_5_6_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_0_ypos.txt",net0.n_5_6_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_0_yneg.txt",net0.n_5_6_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_0_zpos.txt",net0.n_5_6_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_0_zneg.txt",net0.n_5_6_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_1_local.txt",net0.n_5_6_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_1_xpos.txt",net0.n_5_6_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_1_xneg.txt",net0.n_5_6_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_1_ypos.txt",net0.n_5_6_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_1_yneg.txt",net0.n_5_6_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_1_zpos.txt",net0.n_5_6_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_1_zneg.txt",net0.n_5_6_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_1_xpos.txt",net0.n_5_6_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_1_xneg.txt",net0.n_5_6_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_1_ypos.txt",net0.n_5_6_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_1_yneg.txt",net0.n_5_6_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_1_zpos.txt",net0.n_5_6_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_1_zneg.txt",net0.n_5_6_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_1_xpos.txt",net0.n_5_6_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_1_xneg.txt",net0.n_5_6_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_1_ypos.txt",net0.n_5_6_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_1_yneg.txt",net0.n_5_6_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_1_zpos.txt",net0.n_5_6_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_1_zneg.txt",net0.n_5_6_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_2_local.txt",net0.n_5_6_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_2_xpos.txt",net0.n_5_6_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_2_xneg.txt",net0.n_5_6_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_2_ypos.txt",net0.n_5_6_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_2_yneg.txt",net0.n_5_6_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_2_zpos.txt",net0.n_5_6_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_2_zneg.txt",net0.n_5_6_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_2_xpos.txt",net0.n_5_6_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_2_xneg.txt",net0.n_5_6_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_2_ypos.txt",net0.n_5_6_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_2_yneg.txt",net0.n_5_6_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_2_zpos.txt",net0.n_5_6_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_2_zneg.txt",net0.n_5_6_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_2_xpos.txt",net0.n_5_6_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_2_xneg.txt",net0.n_5_6_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_2_ypos.txt",net0.n_5_6_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_2_yneg.txt",net0.n_5_6_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_2_zpos.txt",net0.n_5_6_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_2_zneg.txt",net0.n_5_6_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_3_local.txt",net0.n_5_6_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_3_xpos.txt",net0.n_5_6_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_3_xneg.txt",net0.n_5_6_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_3_ypos.txt",net0.n_5_6_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_3_yneg.txt",net0.n_5_6_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_3_zpos.txt",net0.n_5_6_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_3_zneg.txt",net0.n_5_6_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_3_xpos.txt",net0.n_5_6_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_3_xneg.txt",net0.n_5_6_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_3_ypos.txt",net0.n_5_6_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_3_yneg.txt",net0.n_5_6_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_3_zpos.txt",net0.n_5_6_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_3_zneg.txt",net0.n_5_6_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_3_xpos.txt",net0.n_5_6_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_3_xneg.txt",net0.n_5_6_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_3_ypos.txt",net0.n_5_6_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_3_yneg.txt",net0.n_5_6_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_3_zpos.txt",net0.n_5_6_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_3_zneg.txt",net0.n_5_6_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_4_local.txt",net0.n_5_6_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_4_xpos.txt",net0.n_5_6_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_4_xneg.txt",net0.n_5_6_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_4_ypos.txt",net0.n_5_6_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_4_yneg.txt",net0.n_5_6_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_4_zpos.txt",net0.n_5_6_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_4_zneg.txt",net0.n_5_6_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_4_xpos.txt",net0.n_5_6_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_4_xneg.txt",net0.n_5_6_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_4_ypos.txt",net0.n_5_6_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_4_yneg.txt",net0.n_5_6_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_4_zpos.txt",net0.n_5_6_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_4_zneg.txt",net0.n_5_6_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_4_xpos.txt",net0.n_5_6_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_4_xneg.txt",net0.n_5_6_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_4_ypos.txt",net0.n_5_6_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_4_yneg.txt",net0.n_5_6_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_4_zpos.txt",net0.n_5_6_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_4_zneg.txt",net0.n_5_6_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_5_local.txt",net0.n_5_6_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_5_xpos.txt",net0.n_5_6_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_5_xneg.txt",net0.n_5_6_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_5_ypos.txt",net0.n_5_6_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_5_yneg.txt",net0.n_5_6_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_5_zpos.txt",net0.n_5_6_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_5_zneg.txt",net0.n_5_6_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_5_xpos.txt",net0.n_5_6_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_5_xneg.txt",net0.n_5_6_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_5_ypos.txt",net0.n_5_6_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_5_yneg.txt",net0.n_5_6_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_5_zpos.txt",net0.n_5_6_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_5_zneg.txt",net0.n_5_6_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_5_xpos.txt",net0.n_5_6_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_5_xneg.txt",net0.n_5_6_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_5_ypos.txt",net0.n_5_6_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_5_yneg.txt",net0.n_5_6_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_5_zpos.txt",net0.n_5_6_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_5_zneg.txt",net0.n_5_6_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_6_local.txt",net0.n_5_6_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_6_xpos.txt",net0.n_5_6_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_6_xneg.txt",net0.n_5_6_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_6_ypos.txt",net0.n_5_6_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_6_yneg.txt",net0.n_5_6_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_6_zpos.txt",net0.n_5_6_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_6_zneg.txt",net0.n_5_6_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_6_xpos.txt",net0.n_5_6_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_6_xneg.txt",net0.n_5_6_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_6_ypos.txt",net0.n_5_6_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_6_yneg.txt",net0.n_5_6_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_6_zpos.txt",net0.n_5_6_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_6_zneg.txt",net0.n_5_6_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_6_xpos.txt",net0.n_5_6_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_6_xneg.txt",net0.n_5_6_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_6_ypos.txt",net0.n_5_6_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_6_yneg.txt",net0.n_5_6_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_6_zpos.txt",net0.n_5_6_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_6_zneg.txt",net0.n_5_6_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_7_local.txt",net0.n_5_6_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_7_xpos.txt",net0.n_5_6_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_7_xneg.txt",net0.n_5_6_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_7_ypos.txt",net0.n_5_6_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_7_yneg.txt",net0.n_5_6_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_7_zpos.txt",net0.n_5_6_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_6_7_zneg.txt",net0.n_5_6_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_7_xpos.txt",net0.n_5_6_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_7_xneg.txt",net0.n_5_6_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_7_ypos.txt",net0.n_5_6_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_7_yneg.txt",net0.n_5_6_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_7_zpos.txt",net0.n_5_6_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_6_7_zneg.txt",net0.n_5_6_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_7_xpos.txt",net0.n_5_6_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_7_xneg.txt",net0.n_5_6_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_7_ypos.txt",net0.n_5_6_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_7_yneg.txt",net0.n_5_6_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_7_zpos.txt",net0.n_5_6_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_6_7_zneg.txt",net0.n_5_6_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_0_local.txt",net0.n_5_7_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_0_xpos.txt",net0.n_5_7_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_0_xneg.txt",net0.n_5_7_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_0_ypos.txt",net0.n_5_7_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_0_yneg.txt",net0.n_5_7_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_0_zpos.txt",net0.n_5_7_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_0_zneg.txt",net0.n_5_7_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_0_xpos.txt",net0.n_5_7_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_0_xneg.txt",net0.n_5_7_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_0_ypos.txt",net0.n_5_7_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_0_yneg.txt",net0.n_5_7_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_0_zpos.txt",net0.n_5_7_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_0_zneg.txt",net0.n_5_7_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_0_xpos.txt",net0.n_5_7_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_0_xneg.txt",net0.n_5_7_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_0_ypos.txt",net0.n_5_7_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_0_yneg.txt",net0.n_5_7_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_0_zpos.txt",net0.n_5_7_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_0_zneg.txt",net0.n_5_7_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_1_local.txt",net0.n_5_7_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_1_xpos.txt",net0.n_5_7_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_1_xneg.txt",net0.n_5_7_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_1_ypos.txt",net0.n_5_7_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_1_yneg.txt",net0.n_5_7_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_1_zpos.txt",net0.n_5_7_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_1_zneg.txt",net0.n_5_7_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_1_xpos.txt",net0.n_5_7_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_1_xneg.txt",net0.n_5_7_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_1_ypos.txt",net0.n_5_7_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_1_yneg.txt",net0.n_5_7_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_1_zpos.txt",net0.n_5_7_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_1_zneg.txt",net0.n_5_7_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_1_xpos.txt",net0.n_5_7_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_1_xneg.txt",net0.n_5_7_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_1_ypos.txt",net0.n_5_7_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_1_yneg.txt",net0.n_5_7_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_1_zpos.txt",net0.n_5_7_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_1_zneg.txt",net0.n_5_7_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_2_local.txt",net0.n_5_7_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_2_xpos.txt",net0.n_5_7_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_2_xneg.txt",net0.n_5_7_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_2_ypos.txt",net0.n_5_7_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_2_yneg.txt",net0.n_5_7_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_2_zpos.txt",net0.n_5_7_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_2_zneg.txt",net0.n_5_7_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_2_xpos.txt",net0.n_5_7_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_2_xneg.txt",net0.n_5_7_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_2_ypos.txt",net0.n_5_7_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_2_yneg.txt",net0.n_5_7_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_2_zpos.txt",net0.n_5_7_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_2_zneg.txt",net0.n_5_7_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_2_xpos.txt",net0.n_5_7_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_2_xneg.txt",net0.n_5_7_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_2_ypos.txt",net0.n_5_7_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_2_yneg.txt",net0.n_5_7_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_2_zpos.txt",net0.n_5_7_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_2_zneg.txt",net0.n_5_7_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_3_local.txt",net0.n_5_7_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_3_xpos.txt",net0.n_5_7_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_3_xneg.txt",net0.n_5_7_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_3_ypos.txt",net0.n_5_7_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_3_yneg.txt",net0.n_5_7_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_3_zpos.txt",net0.n_5_7_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_3_zneg.txt",net0.n_5_7_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_3_xpos.txt",net0.n_5_7_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_3_xneg.txt",net0.n_5_7_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_3_ypos.txt",net0.n_5_7_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_3_yneg.txt",net0.n_5_7_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_3_zpos.txt",net0.n_5_7_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_3_zneg.txt",net0.n_5_7_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_3_xpos.txt",net0.n_5_7_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_3_xneg.txt",net0.n_5_7_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_3_ypos.txt",net0.n_5_7_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_3_yneg.txt",net0.n_5_7_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_3_zpos.txt",net0.n_5_7_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_3_zneg.txt",net0.n_5_7_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_4_local.txt",net0.n_5_7_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_4_xpos.txt",net0.n_5_7_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_4_xneg.txt",net0.n_5_7_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_4_ypos.txt",net0.n_5_7_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_4_yneg.txt",net0.n_5_7_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_4_zpos.txt",net0.n_5_7_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_4_zneg.txt",net0.n_5_7_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_4_xpos.txt",net0.n_5_7_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_4_xneg.txt",net0.n_5_7_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_4_ypos.txt",net0.n_5_7_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_4_yneg.txt",net0.n_5_7_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_4_zpos.txt",net0.n_5_7_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_4_zneg.txt",net0.n_5_7_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_4_xpos.txt",net0.n_5_7_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_4_xneg.txt",net0.n_5_7_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_4_ypos.txt",net0.n_5_7_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_4_yneg.txt",net0.n_5_7_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_4_zpos.txt",net0.n_5_7_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_4_zneg.txt",net0.n_5_7_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_5_local.txt",net0.n_5_7_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_5_xpos.txt",net0.n_5_7_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_5_xneg.txt",net0.n_5_7_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_5_ypos.txt",net0.n_5_7_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_5_yneg.txt",net0.n_5_7_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_5_zpos.txt",net0.n_5_7_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_5_zneg.txt",net0.n_5_7_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_5_xpos.txt",net0.n_5_7_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_5_xneg.txt",net0.n_5_7_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_5_ypos.txt",net0.n_5_7_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_5_yneg.txt",net0.n_5_7_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_5_zpos.txt",net0.n_5_7_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_5_zneg.txt",net0.n_5_7_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_5_xpos.txt",net0.n_5_7_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_5_xneg.txt",net0.n_5_7_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_5_ypos.txt",net0.n_5_7_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_5_yneg.txt",net0.n_5_7_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_5_zpos.txt",net0.n_5_7_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_5_zneg.txt",net0.n_5_7_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_6_local.txt",net0.n_5_7_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_6_xpos.txt",net0.n_5_7_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_6_xneg.txt",net0.n_5_7_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_6_ypos.txt",net0.n_5_7_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_6_yneg.txt",net0.n_5_7_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_6_zpos.txt",net0.n_5_7_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_6_zneg.txt",net0.n_5_7_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_6_xpos.txt",net0.n_5_7_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_6_xneg.txt",net0.n_5_7_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_6_ypos.txt",net0.n_5_7_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_6_yneg.txt",net0.n_5_7_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_6_zpos.txt",net0.n_5_7_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_6_zneg.txt",net0.n_5_7_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_6_xpos.txt",net0.n_5_7_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_6_xneg.txt",net0.n_5_7_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_6_ypos.txt",net0.n_5_7_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_6_yneg.txt",net0.n_5_7_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_6_zpos.txt",net0.n_5_7_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_6_zneg.txt",net0.n_5_7_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_7_local.txt",net0.n_5_7_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_7_xpos.txt",net0.n_5_7_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_7_xneg.txt",net0.n_5_7_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_7_ypos.txt",net0.n_5_7_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_7_yneg.txt",net0.n_5_7_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_7_zpos.txt",net0.n_5_7_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_5_7_7_zneg.txt",net0.n_5_7_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_7_xpos.txt",net0.n_5_7_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_7_xneg.txt",net0.n_5_7_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_7_ypos.txt",net0.n_5_7_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_7_yneg.txt",net0.n_5_7_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_7_zpos.txt",net0.n_5_7_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_5_7_7_zneg.txt",net0.n_5_7_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_7_xpos.txt",net0.n_5_7_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_7_xneg.txt",net0.n_5_7_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_7_ypos.txt",net0.n_5_7_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_7_yneg.txt",net0.n_5_7_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_7_zpos.txt",net0.n_5_7_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_5_7_7_zneg.txt",net0.n_5_7_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_0_local.txt",net0.n_6_0_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_0_xpos.txt",net0.n_6_0_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_0_xneg.txt",net0.n_6_0_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_0_ypos.txt",net0.n_6_0_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_0_yneg.txt",net0.n_6_0_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_0_zpos.txt",net0.n_6_0_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_0_zneg.txt",net0.n_6_0_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_0_xpos.txt",net0.n_6_0_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_0_xneg.txt",net0.n_6_0_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_0_ypos.txt",net0.n_6_0_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_0_yneg.txt",net0.n_6_0_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_0_zpos.txt",net0.n_6_0_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_0_zneg.txt",net0.n_6_0_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_0_xpos.txt",net0.n_6_0_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_0_xneg.txt",net0.n_6_0_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_0_ypos.txt",net0.n_6_0_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_0_yneg.txt",net0.n_6_0_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_0_zpos.txt",net0.n_6_0_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_0_zneg.txt",net0.n_6_0_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_1_local.txt",net0.n_6_0_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_1_xpos.txt",net0.n_6_0_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_1_xneg.txt",net0.n_6_0_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_1_ypos.txt",net0.n_6_0_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_1_yneg.txt",net0.n_6_0_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_1_zpos.txt",net0.n_6_0_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_1_zneg.txt",net0.n_6_0_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_1_xpos.txt",net0.n_6_0_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_1_xneg.txt",net0.n_6_0_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_1_ypos.txt",net0.n_6_0_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_1_yneg.txt",net0.n_6_0_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_1_zpos.txt",net0.n_6_0_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_1_zneg.txt",net0.n_6_0_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_1_xpos.txt",net0.n_6_0_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_1_xneg.txt",net0.n_6_0_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_1_ypos.txt",net0.n_6_0_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_1_yneg.txt",net0.n_6_0_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_1_zpos.txt",net0.n_6_0_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_1_zneg.txt",net0.n_6_0_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_2_local.txt",net0.n_6_0_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_2_xpos.txt",net0.n_6_0_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_2_xneg.txt",net0.n_6_0_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_2_ypos.txt",net0.n_6_0_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_2_yneg.txt",net0.n_6_0_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_2_zpos.txt",net0.n_6_0_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_2_zneg.txt",net0.n_6_0_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_2_xpos.txt",net0.n_6_0_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_2_xneg.txt",net0.n_6_0_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_2_ypos.txt",net0.n_6_0_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_2_yneg.txt",net0.n_6_0_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_2_zpos.txt",net0.n_6_0_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_2_zneg.txt",net0.n_6_0_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_2_xpos.txt",net0.n_6_0_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_2_xneg.txt",net0.n_6_0_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_2_ypos.txt",net0.n_6_0_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_2_yneg.txt",net0.n_6_0_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_2_zpos.txt",net0.n_6_0_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_2_zneg.txt",net0.n_6_0_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_3_local.txt",net0.n_6_0_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_3_xpos.txt",net0.n_6_0_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_3_xneg.txt",net0.n_6_0_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_3_ypos.txt",net0.n_6_0_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_3_yneg.txt",net0.n_6_0_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_3_zpos.txt",net0.n_6_0_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_3_zneg.txt",net0.n_6_0_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_3_xpos.txt",net0.n_6_0_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_3_xneg.txt",net0.n_6_0_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_3_ypos.txt",net0.n_6_0_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_3_yneg.txt",net0.n_6_0_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_3_zpos.txt",net0.n_6_0_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_3_zneg.txt",net0.n_6_0_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_3_xpos.txt",net0.n_6_0_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_3_xneg.txt",net0.n_6_0_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_3_ypos.txt",net0.n_6_0_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_3_yneg.txt",net0.n_6_0_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_3_zpos.txt",net0.n_6_0_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_3_zneg.txt",net0.n_6_0_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_4_local.txt",net0.n_6_0_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_4_xpos.txt",net0.n_6_0_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_4_xneg.txt",net0.n_6_0_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_4_ypos.txt",net0.n_6_0_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_4_yneg.txt",net0.n_6_0_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_4_zpos.txt",net0.n_6_0_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_4_zneg.txt",net0.n_6_0_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_4_xpos.txt",net0.n_6_0_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_4_xneg.txt",net0.n_6_0_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_4_ypos.txt",net0.n_6_0_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_4_yneg.txt",net0.n_6_0_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_4_zpos.txt",net0.n_6_0_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_4_zneg.txt",net0.n_6_0_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_4_xpos.txt",net0.n_6_0_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_4_xneg.txt",net0.n_6_0_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_4_ypos.txt",net0.n_6_0_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_4_yneg.txt",net0.n_6_0_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_4_zpos.txt",net0.n_6_0_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_4_zneg.txt",net0.n_6_0_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_5_local.txt",net0.n_6_0_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_5_xpos.txt",net0.n_6_0_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_5_xneg.txt",net0.n_6_0_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_5_ypos.txt",net0.n_6_0_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_5_yneg.txt",net0.n_6_0_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_5_zpos.txt",net0.n_6_0_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_5_zneg.txt",net0.n_6_0_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_5_xpos.txt",net0.n_6_0_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_5_xneg.txt",net0.n_6_0_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_5_ypos.txt",net0.n_6_0_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_5_yneg.txt",net0.n_6_0_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_5_zpos.txt",net0.n_6_0_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_5_zneg.txt",net0.n_6_0_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_5_xpos.txt",net0.n_6_0_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_5_xneg.txt",net0.n_6_0_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_5_ypos.txt",net0.n_6_0_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_5_yneg.txt",net0.n_6_0_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_5_zpos.txt",net0.n_6_0_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_5_zneg.txt",net0.n_6_0_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_6_local.txt",net0.n_6_0_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_6_xpos.txt",net0.n_6_0_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_6_xneg.txt",net0.n_6_0_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_6_ypos.txt",net0.n_6_0_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_6_yneg.txt",net0.n_6_0_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_6_zpos.txt",net0.n_6_0_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_6_zneg.txt",net0.n_6_0_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_6_xpos.txt",net0.n_6_0_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_6_xneg.txt",net0.n_6_0_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_6_ypos.txt",net0.n_6_0_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_6_yneg.txt",net0.n_6_0_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_6_zpos.txt",net0.n_6_0_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_6_zneg.txt",net0.n_6_0_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_6_xpos.txt",net0.n_6_0_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_6_xneg.txt",net0.n_6_0_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_6_ypos.txt",net0.n_6_0_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_6_yneg.txt",net0.n_6_0_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_6_zpos.txt",net0.n_6_0_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_6_zneg.txt",net0.n_6_0_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_7_local.txt",net0.n_6_0_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_7_xpos.txt",net0.n_6_0_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_7_xneg.txt",net0.n_6_0_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_7_ypos.txt",net0.n_6_0_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_7_yneg.txt",net0.n_6_0_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_7_zpos.txt",net0.n_6_0_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_0_7_zneg.txt",net0.n_6_0_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_7_xpos.txt",net0.n_6_0_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_7_xneg.txt",net0.n_6_0_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_7_ypos.txt",net0.n_6_0_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_7_yneg.txt",net0.n_6_0_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_7_zpos.txt",net0.n_6_0_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_0_7_zneg.txt",net0.n_6_0_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_7_xpos.txt",net0.n_6_0_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_7_xneg.txt",net0.n_6_0_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_7_ypos.txt",net0.n_6_0_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_7_yneg.txt",net0.n_6_0_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_7_zpos.txt",net0.n_6_0_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_0_7_zneg.txt",net0.n_6_0_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_0_local.txt",net0.n_6_1_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_0_xpos.txt",net0.n_6_1_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_0_xneg.txt",net0.n_6_1_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_0_ypos.txt",net0.n_6_1_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_0_yneg.txt",net0.n_6_1_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_0_zpos.txt",net0.n_6_1_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_0_zneg.txt",net0.n_6_1_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_0_xpos.txt",net0.n_6_1_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_0_xneg.txt",net0.n_6_1_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_0_ypos.txt",net0.n_6_1_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_0_yneg.txt",net0.n_6_1_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_0_zpos.txt",net0.n_6_1_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_0_zneg.txt",net0.n_6_1_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_0_xpos.txt",net0.n_6_1_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_0_xneg.txt",net0.n_6_1_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_0_ypos.txt",net0.n_6_1_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_0_yneg.txt",net0.n_6_1_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_0_zpos.txt",net0.n_6_1_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_0_zneg.txt",net0.n_6_1_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_1_local.txt",net0.n_6_1_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_1_xpos.txt",net0.n_6_1_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_1_xneg.txt",net0.n_6_1_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_1_ypos.txt",net0.n_6_1_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_1_yneg.txt",net0.n_6_1_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_1_zpos.txt",net0.n_6_1_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_1_zneg.txt",net0.n_6_1_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_1_xpos.txt",net0.n_6_1_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_1_xneg.txt",net0.n_6_1_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_1_ypos.txt",net0.n_6_1_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_1_yneg.txt",net0.n_6_1_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_1_zpos.txt",net0.n_6_1_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_1_zneg.txt",net0.n_6_1_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_1_xpos.txt",net0.n_6_1_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_1_xneg.txt",net0.n_6_1_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_1_ypos.txt",net0.n_6_1_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_1_yneg.txt",net0.n_6_1_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_1_zpos.txt",net0.n_6_1_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_1_zneg.txt",net0.n_6_1_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_2_local.txt",net0.n_6_1_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_2_xpos.txt",net0.n_6_1_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_2_xneg.txt",net0.n_6_1_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_2_ypos.txt",net0.n_6_1_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_2_yneg.txt",net0.n_6_1_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_2_zpos.txt",net0.n_6_1_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_2_zneg.txt",net0.n_6_1_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_2_xpos.txt",net0.n_6_1_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_2_xneg.txt",net0.n_6_1_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_2_ypos.txt",net0.n_6_1_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_2_yneg.txt",net0.n_6_1_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_2_zpos.txt",net0.n_6_1_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_2_zneg.txt",net0.n_6_1_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_2_xpos.txt",net0.n_6_1_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_2_xneg.txt",net0.n_6_1_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_2_ypos.txt",net0.n_6_1_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_2_yneg.txt",net0.n_6_1_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_2_zpos.txt",net0.n_6_1_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_2_zneg.txt",net0.n_6_1_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_3_local.txt",net0.n_6_1_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_3_xpos.txt",net0.n_6_1_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_3_xneg.txt",net0.n_6_1_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_3_ypos.txt",net0.n_6_1_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_3_yneg.txt",net0.n_6_1_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_3_zpos.txt",net0.n_6_1_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_3_zneg.txt",net0.n_6_1_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_3_xpos.txt",net0.n_6_1_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_3_xneg.txt",net0.n_6_1_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_3_ypos.txt",net0.n_6_1_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_3_yneg.txt",net0.n_6_1_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_3_zpos.txt",net0.n_6_1_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_3_zneg.txt",net0.n_6_1_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_3_xpos.txt",net0.n_6_1_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_3_xneg.txt",net0.n_6_1_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_3_ypos.txt",net0.n_6_1_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_3_yneg.txt",net0.n_6_1_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_3_zpos.txt",net0.n_6_1_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_3_zneg.txt",net0.n_6_1_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_4_local.txt",net0.n_6_1_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_4_xpos.txt",net0.n_6_1_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_4_xneg.txt",net0.n_6_1_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_4_ypos.txt",net0.n_6_1_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_4_yneg.txt",net0.n_6_1_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_4_zpos.txt",net0.n_6_1_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_4_zneg.txt",net0.n_6_1_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_4_xpos.txt",net0.n_6_1_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_4_xneg.txt",net0.n_6_1_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_4_ypos.txt",net0.n_6_1_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_4_yneg.txt",net0.n_6_1_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_4_zpos.txt",net0.n_6_1_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_4_zneg.txt",net0.n_6_1_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_4_xpos.txt",net0.n_6_1_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_4_xneg.txt",net0.n_6_1_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_4_ypos.txt",net0.n_6_1_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_4_yneg.txt",net0.n_6_1_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_4_zpos.txt",net0.n_6_1_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_4_zneg.txt",net0.n_6_1_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_5_local.txt",net0.n_6_1_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_5_xpos.txt",net0.n_6_1_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_5_xneg.txt",net0.n_6_1_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_5_ypos.txt",net0.n_6_1_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_5_yneg.txt",net0.n_6_1_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_5_zpos.txt",net0.n_6_1_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_5_zneg.txt",net0.n_6_1_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_5_xpos.txt",net0.n_6_1_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_5_xneg.txt",net0.n_6_1_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_5_ypos.txt",net0.n_6_1_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_5_yneg.txt",net0.n_6_1_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_5_zpos.txt",net0.n_6_1_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_5_zneg.txt",net0.n_6_1_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_5_xpos.txt",net0.n_6_1_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_5_xneg.txt",net0.n_6_1_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_5_ypos.txt",net0.n_6_1_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_5_yneg.txt",net0.n_6_1_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_5_zpos.txt",net0.n_6_1_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_5_zneg.txt",net0.n_6_1_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_6_local.txt",net0.n_6_1_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_6_xpos.txt",net0.n_6_1_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_6_xneg.txt",net0.n_6_1_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_6_ypos.txt",net0.n_6_1_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_6_yneg.txt",net0.n_6_1_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_6_zpos.txt",net0.n_6_1_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_6_zneg.txt",net0.n_6_1_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_6_xpos.txt",net0.n_6_1_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_6_xneg.txt",net0.n_6_1_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_6_ypos.txt",net0.n_6_1_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_6_yneg.txt",net0.n_6_1_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_6_zpos.txt",net0.n_6_1_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_6_zneg.txt",net0.n_6_1_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_6_xpos.txt",net0.n_6_1_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_6_xneg.txt",net0.n_6_1_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_6_ypos.txt",net0.n_6_1_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_6_yneg.txt",net0.n_6_1_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_6_zpos.txt",net0.n_6_1_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_6_zneg.txt",net0.n_6_1_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_7_local.txt",net0.n_6_1_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_7_xpos.txt",net0.n_6_1_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_7_xneg.txt",net0.n_6_1_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_7_ypos.txt",net0.n_6_1_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_7_yneg.txt",net0.n_6_1_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_7_zpos.txt",net0.n_6_1_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_1_7_zneg.txt",net0.n_6_1_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_7_xpos.txt",net0.n_6_1_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_7_xneg.txt",net0.n_6_1_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_7_ypos.txt",net0.n_6_1_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_7_yneg.txt",net0.n_6_1_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_7_zpos.txt",net0.n_6_1_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_1_7_zneg.txt",net0.n_6_1_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_7_xpos.txt",net0.n_6_1_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_7_xneg.txt",net0.n_6_1_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_7_ypos.txt",net0.n_6_1_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_7_yneg.txt",net0.n_6_1_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_7_zpos.txt",net0.n_6_1_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_1_7_zneg.txt",net0.n_6_1_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_0_local.txt",net0.n_6_2_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_0_xpos.txt",net0.n_6_2_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_0_xneg.txt",net0.n_6_2_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_0_ypos.txt",net0.n_6_2_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_0_yneg.txt",net0.n_6_2_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_0_zpos.txt",net0.n_6_2_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_0_zneg.txt",net0.n_6_2_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_0_xpos.txt",net0.n_6_2_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_0_xneg.txt",net0.n_6_2_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_0_ypos.txt",net0.n_6_2_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_0_yneg.txt",net0.n_6_2_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_0_zpos.txt",net0.n_6_2_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_0_zneg.txt",net0.n_6_2_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_0_xpos.txt",net0.n_6_2_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_0_xneg.txt",net0.n_6_2_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_0_ypos.txt",net0.n_6_2_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_0_yneg.txt",net0.n_6_2_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_0_zpos.txt",net0.n_6_2_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_0_zneg.txt",net0.n_6_2_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_1_local.txt",net0.n_6_2_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_1_xpos.txt",net0.n_6_2_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_1_xneg.txt",net0.n_6_2_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_1_ypos.txt",net0.n_6_2_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_1_yneg.txt",net0.n_6_2_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_1_zpos.txt",net0.n_6_2_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_1_zneg.txt",net0.n_6_2_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_1_xpos.txt",net0.n_6_2_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_1_xneg.txt",net0.n_6_2_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_1_ypos.txt",net0.n_6_2_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_1_yneg.txt",net0.n_6_2_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_1_zpos.txt",net0.n_6_2_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_1_zneg.txt",net0.n_6_2_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_1_xpos.txt",net0.n_6_2_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_1_xneg.txt",net0.n_6_2_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_1_ypos.txt",net0.n_6_2_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_1_yneg.txt",net0.n_6_2_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_1_zpos.txt",net0.n_6_2_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_1_zneg.txt",net0.n_6_2_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_2_local.txt",net0.n_6_2_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_2_xpos.txt",net0.n_6_2_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_2_xneg.txt",net0.n_6_2_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_2_ypos.txt",net0.n_6_2_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_2_yneg.txt",net0.n_6_2_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_2_zpos.txt",net0.n_6_2_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_2_zneg.txt",net0.n_6_2_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_2_xpos.txt",net0.n_6_2_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_2_xneg.txt",net0.n_6_2_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_2_ypos.txt",net0.n_6_2_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_2_yneg.txt",net0.n_6_2_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_2_zpos.txt",net0.n_6_2_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_2_zneg.txt",net0.n_6_2_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_2_xpos.txt",net0.n_6_2_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_2_xneg.txt",net0.n_6_2_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_2_ypos.txt",net0.n_6_2_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_2_yneg.txt",net0.n_6_2_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_2_zpos.txt",net0.n_6_2_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_2_zneg.txt",net0.n_6_2_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_3_local.txt",net0.n_6_2_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_3_xpos.txt",net0.n_6_2_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_3_xneg.txt",net0.n_6_2_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_3_ypos.txt",net0.n_6_2_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_3_yneg.txt",net0.n_6_2_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_3_zpos.txt",net0.n_6_2_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_3_zneg.txt",net0.n_6_2_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_3_xpos.txt",net0.n_6_2_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_3_xneg.txt",net0.n_6_2_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_3_ypos.txt",net0.n_6_2_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_3_yneg.txt",net0.n_6_2_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_3_zpos.txt",net0.n_6_2_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_3_zneg.txt",net0.n_6_2_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_3_xpos.txt",net0.n_6_2_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_3_xneg.txt",net0.n_6_2_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_3_ypos.txt",net0.n_6_2_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_3_yneg.txt",net0.n_6_2_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_3_zpos.txt",net0.n_6_2_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_3_zneg.txt",net0.n_6_2_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_4_local.txt",net0.n_6_2_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_4_xpos.txt",net0.n_6_2_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_4_xneg.txt",net0.n_6_2_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_4_ypos.txt",net0.n_6_2_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_4_yneg.txt",net0.n_6_2_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_4_zpos.txt",net0.n_6_2_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_4_zneg.txt",net0.n_6_2_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_4_xpos.txt",net0.n_6_2_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_4_xneg.txt",net0.n_6_2_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_4_ypos.txt",net0.n_6_2_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_4_yneg.txt",net0.n_6_2_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_4_zpos.txt",net0.n_6_2_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_4_zneg.txt",net0.n_6_2_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_4_xpos.txt",net0.n_6_2_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_4_xneg.txt",net0.n_6_2_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_4_ypos.txt",net0.n_6_2_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_4_yneg.txt",net0.n_6_2_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_4_zpos.txt",net0.n_6_2_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_4_zneg.txt",net0.n_6_2_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_5_local.txt",net0.n_6_2_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_5_xpos.txt",net0.n_6_2_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_5_xneg.txt",net0.n_6_2_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_5_ypos.txt",net0.n_6_2_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_5_yneg.txt",net0.n_6_2_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_5_zpos.txt",net0.n_6_2_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_5_zneg.txt",net0.n_6_2_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_5_xpos.txt",net0.n_6_2_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_5_xneg.txt",net0.n_6_2_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_5_ypos.txt",net0.n_6_2_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_5_yneg.txt",net0.n_6_2_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_5_zpos.txt",net0.n_6_2_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_5_zneg.txt",net0.n_6_2_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_5_xpos.txt",net0.n_6_2_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_5_xneg.txt",net0.n_6_2_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_5_ypos.txt",net0.n_6_2_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_5_yneg.txt",net0.n_6_2_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_5_zpos.txt",net0.n_6_2_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_5_zneg.txt",net0.n_6_2_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_6_local.txt",net0.n_6_2_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_6_xpos.txt",net0.n_6_2_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_6_xneg.txt",net0.n_6_2_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_6_ypos.txt",net0.n_6_2_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_6_yneg.txt",net0.n_6_2_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_6_zpos.txt",net0.n_6_2_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_6_zneg.txt",net0.n_6_2_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_6_xpos.txt",net0.n_6_2_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_6_xneg.txt",net0.n_6_2_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_6_ypos.txt",net0.n_6_2_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_6_yneg.txt",net0.n_6_2_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_6_zpos.txt",net0.n_6_2_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_6_zneg.txt",net0.n_6_2_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_6_xpos.txt",net0.n_6_2_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_6_xneg.txt",net0.n_6_2_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_6_ypos.txt",net0.n_6_2_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_6_yneg.txt",net0.n_6_2_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_6_zpos.txt",net0.n_6_2_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_6_zneg.txt",net0.n_6_2_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_7_local.txt",net0.n_6_2_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_7_xpos.txt",net0.n_6_2_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_7_xneg.txt",net0.n_6_2_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_7_ypos.txt",net0.n_6_2_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_7_yneg.txt",net0.n_6_2_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_7_zpos.txt",net0.n_6_2_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_2_7_zneg.txt",net0.n_6_2_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_7_xpos.txt",net0.n_6_2_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_7_xneg.txt",net0.n_6_2_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_7_ypos.txt",net0.n_6_2_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_7_yneg.txt",net0.n_6_2_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_7_zpos.txt",net0.n_6_2_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_2_7_zneg.txt",net0.n_6_2_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_7_xpos.txt",net0.n_6_2_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_7_xneg.txt",net0.n_6_2_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_7_ypos.txt",net0.n_6_2_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_7_yneg.txt",net0.n_6_2_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_7_zpos.txt",net0.n_6_2_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_2_7_zneg.txt",net0.n_6_2_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_0_local.txt",net0.n_6_3_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_0_xpos.txt",net0.n_6_3_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_0_xneg.txt",net0.n_6_3_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_0_ypos.txt",net0.n_6_3_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_0_yneg.txt",net0.n_6_3_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_0_zpos.txt",net0.n_6_3_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_0_zneg.txt",net0.n_6_3_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_0_xpos.txt",net0.n_6_3_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_0_xneg.txt",net0.n_6_3_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_0_ypos.txt",net0.n_6_3_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_0_yneg.txt",net0.n_6_3_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_0_zpos.txt",net0.n_6_3_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_0_zneg.txt",net0.n_6_3_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_0_xpos.txt",net0.n_6_3_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_0_xneg.txt",net0.n_6_3_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_0_ypos.txt",net0.n_6_3_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_0_yneg.txt",net0.n_6_3_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_0_zpos.txt",net0.n_6_3_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_0_zneg.txt",net0.n_6_3_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_1_local.txt",net0.n_6_3_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_1_xpos.txt",net0.n_6_3_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_1_xneg.txt",net0.n_6_3_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_1_ypos.txt",net0.n_6_3_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_1_yneg.txt",net0.n_6_3_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_1_zpos.txt",net0.n_6_3_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_1_zneg.txt",net0.n_6_3_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_1_xpos.txt",net0.n_6_3_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_1_xneg.txt",net0.n_6_3_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_1_ypos.txt",net0.n_6_3_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_1_yneg.txt",net0.n_6_3_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_1_zpos.txt",net0.n_6_3_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_1_zneg.txt",net0.n_6_3_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_1_xpos.txt",net0.n_6_3_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_1_xneg.txt",net0.n_6_3_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_1_ypos.txt",net0.n_6_3_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_1_yneg.txt",net0.n_6_3_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_1_zpos.txt",net0.n_6_3_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_1_zneg.txt",net0.n_6_3_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_2_local.txt",net0.n_6_3_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_2_xpos.txt",net0.n_6_3_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_2_xneg.txt",net0.n_6_3_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_2_ypos.txt",net0.n_6_3_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_2_yneg.txt",net0.n_6_3_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_2_zpos.txt",net0.n_6_3_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_2_zneg.txt",net0.n_6_3_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_2_xpos.txt",net0.n_6_3_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_2_xneg.txt",net0.n_6_3_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_2_ypos.txt",net0.n_6_3_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_2_yneg.txt",net0.n_6_3_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_2_zpos.txt",net0.n_6_3_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_2_zneg.txt",net0.n_6_3_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_2_xpos.txt",net0.n_6_3_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_2_xneg.txt",net0.n_6_3_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_2_ypos.txt",net0.n_6_3_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_2_yneg.txt",net0.n_6_3_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_2_zpos.txt",net0.n_6_3_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_2_zneg.txt",net0.n_6_3_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_3_local.txt",net0.n_6_3_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_3_xpos.txt",net0.n_6_3_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_3_xneg.txt",net0.n_6_3_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_3_ypos.txt",net0.n_6_3_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_3_yneg.txt",net0.n_6_3_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_3_zpos.txt",net0.n_6_3_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_3_zneg.txt",net0.n_6_3_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_3_xpos.txt",net0.n_6_3_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_3_xneg.txt",net0.n_6_3_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_3_ypos.txt",net0.n_6_3_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_3_yneg.txt",net0.n_6_3_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_3_zpos.txt",net0.n_6_3_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_3_zneg.txt",net0.n_6_3_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_3_xpos.txt",net0.n_6_3_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_3_xneg.txt",net0.n_6_3_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_3_ypos.txt",net0.n_6_3_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_3_yneg.txt",net0.n_6_3_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_3_zpos.txt",net0.n_6_3_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_3_zneg.txt",net0.n_6_3_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_4_local.txt",net0.n_6_3_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_4_xpos.txt",net0.n_6_3_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_4_xneg.txt",net0.n_6_3_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_4_ypos.txt",net0.n_6_3_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_4_yneg.txt",net0.n_6_3_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_4_zpos.txt",net0.n_6_3_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_4_zneg.txt",net0.n_6_3_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_4_xpos.txt",net0.n_6_3_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_4_xneg.txt",net0.n_6_3_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_4_ypos.txt",net0.n_6_3_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_4_yneg.txt",net0.n_6_3_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_4_zpos.txt",net0.n_6_3_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_4_zneg.txt",net0.n_6_3_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_4_xpos.txt",net0.n_6_3_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_4_xneg.txt",net0.n_6_3_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_4_ypos.txt",net0.n_6_3_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_4_yneg.txt",net0.n_6_3_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_4_zpos.txt",net0.n_6_3_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_4_zneg.txt",net0.n_6_3_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_5_local.txt",net0.n_6_3_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_5_xpos.txt",net0.n_6_3_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_5_xneg.txt",net0.n_6_3_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_5_ypos.txt",net0.n_6_3_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_5_yneg.txt",net0.n_6_3_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_5_zpos.txt",net0.n_6_3_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_5_zneg.txt",net0.n_6_3_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_5_xpos.txt",net0.n_6_3_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_5_xneg.txt",net0.n_6_3_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_5_ypos.txt",net0.n_6_3_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_5_yneg.txt",net0.n_6_3_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_5_zpos.txt",net0.n_6_3_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_5_zneg.txt",net0.n_6_3_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_5_xpos.txt",net0.n_6_3_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_5_xneg.txt",net0.n_6_3_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_5_ypos.txt",net0.n_6_3_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_5_yneg.txt",net0.n_6_3_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_5_zpos.txt",net0.n_6_3_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_5_zneg.txt",net0.n_6_3_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_6_local.txt",net0.n_6_3_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_6_xpos.txt",net0.n_6_3_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_6_xneg.txt",net0.n_6_3_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_6_ypos.txt",net0.n_6_3_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_6_yneg.txt",net0.n_6_3_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_6_zpos.txt",net0.n_6_3_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_6_zneg.txt",net0.n_6_3_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_6_xpos.txt",net0.n_6_3_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_6_xneg.txt",net0.n_6_3_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_6_ypos.txt",net0.n_6_3_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_6_yneg.txt",net0.n_6_3_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_6_zpos.txt",net0.n_6_3_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_6_zneg.txt",net0.n_6_3_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_6_xpos.txt",net0.n_6_3_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_6_xneg.txt",net0.n_6_3_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_6_ypos.txt",net0.n_6_3_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_6_yneg.txt",net0.n_6_3_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_6_zpos.txt",net0.n_6_3_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_6_zneg.txt",net0.n_6_3_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_7_local.txt",net0.n_6_3_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_7_xpos.txt",net0.n_6_3_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_7_xneg.txt",net0.n_6_3_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_7_ypos.txt",net0.n_6_3_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_7_yneg.txt",net0.n_6_3_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_7_zpos.txt",net0.n_6_3_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_3_7_zneg.txt",net0.n_6_3_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_7_xpos.txt",net0.n_6_3_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_7_xneg.txt",net0.n_6_3_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_7_ypos.txt",net0.n_6_3_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_7_yneg.txt",net0.n_6_3_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_7_zpos.txt",net0.n_6_3_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_3_7_zneg.txt",net0.n_6_3_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_7_xpos.txt",net0.n_6_3_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_7_xneg.txt",net0.n_6_3_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_7_ypos.txt",net0.n_6_3_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_7_yneg.txt",net0.n_6_3_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_7_zpos.txt",net0.n_6_3_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_3_7_zneg.txt",net0.n_6_3_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_0_local.txt",net0.n_6_4_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_0_xpos.txt",net0.n_6_4_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_0_xneg.txt",net0.n_6_4_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_0_ypos.txt",net0.n_6_4_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_0_yneg.txt",net0.n_6_4_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_0_zpos.txt",net0.n_6_4_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_0_zneg.txt",net0.n_6_4_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_0_xpos.txt",net0.n_6_4_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_0_xneg.txt",net0.n_6_4_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_0_ypos.txt",net0.n_6_4_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_0_yneg.txt",net0.n_6_4_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_0_zpos.txt",net0.n_6_4_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_0_zneg.txt",net0.n_6_4_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_0_xpos.txt",net0.n_6_4_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_0_xneg.txt",net0.n_6_4_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_0_ypos.txt",net0.n_6_4_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_0_yneg.txt",net0.n_6_4_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_0_zpos.txt",net0.n_6_4_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_0_zneg.txt",net0.n_6_4_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_1_local.txt",net0.n_6_4_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_1_xpos.txt",net0.n_6_4_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_1_xneg.txt",net0.n_6_4_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_1_ypos.txt",net0.n_6_4_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_1_yneg.txt",net0.n_6_4_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_1_zpos.txt",net0.n_6_4_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_1_zneg.txt",net0.n_6_4_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_1_xpos.txt",net0.n_6_4_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_1_xneg.txt",net0.n_6_4_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_1_ypos.txt",net0.n_6_4_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_1_yneg.txt",net0.n_6_4_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_1_zpos.txt",net0.n_6_4_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_1_zneg.txt",net0.n_6_4_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_1_xpos.txt",net0.n_6_4_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_1_xneg.txt",net0.n_6_4_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_1_ypos.txt",net0.n_6_4_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_1_yneg.txt",net0.n_6_4_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_1_zpos.txt",net0.n_6_4_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_1_zneg.txt",net0.n_6_4_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_2_local.txt",net0.n_6_4_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_2_xpos.txt",net0.n_6_4_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_2_xneg.txt",net0.n_6_4_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_2_ypos.txt",net0.n_6_4_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_2_yneg.txt",net0.n_6_4_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_2_zpos.txt",net0.n_6_4_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_2_zneg.txt",net0.n_6_4_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_2_xpos.txt",net0.n_6_4_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_2_xneg.txt",net0.n_6_4_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_2_ypos.txt",net0.n_6_4_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_2_yneg.txt",net0.n_6_4_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_2_zpos.txt",net0.n_6_4_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_2_zneg.txt",net0.n_6_4_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_2_xpos.txt",net0.n_6_4_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_2_xneg.txt",net0.n_6_4_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_2_ypos.txt",net0.n_6_4_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_2_yneg.txt",net0.n_6_4_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_2_zpos.txt",net0.n_6_4_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_2_zneg.txt",net0.n_6_4_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_3_local.txt",net0.n_6_4_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_3_xpos.txt",net0.n_6_4_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_3_xneg.txt",net0.n_6_4_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_3_ypos.txt",net0.n_6_4_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_3_yneg.txt",net0.n_6_4_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_3_zpos.txt",net0.n_6_4_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_3_zneg.txt",net0.n_6_4_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_3_xpos.txt",net0.n_6_4_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_3_xneg.txt",net0.n_6_4_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_3_ypos.txt",net0.n_6_4_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_3_yneg.txt",net0.n_6_4_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_3_zpos.txt",net0.n_6_4_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_3_zneg.txt",net0.n_6_4_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_3_xpos.txt",net0.n_6_4_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_3_xneg.txt",net0.n_6_4_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_3_ypos.txt",net0.n_6_4_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_3_yneg.txt",net0.n_6_4_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_3_zpos.txt",net0.n_6_4_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_3_zneg.txt",net0.n_6_4_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_4_local.txt",net0.n_6_4_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_4_xpos.txt",net0.n_6_4_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_4_xneg.txt",net0.n_6_4_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_4_ypos.txt",net0.n_6_4_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_4_yneg.txt",net0.n_6_4_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_4_zpos.txt",net0.n_6_4_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_4_zneg.txt",net0.n_6_4_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_4_xpos.txt",net0.n_6_4_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_4_xneg.txt",net0.n_6_4_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_4_ypos.txt",net0.n_6_4_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_4_yneg.txt",net0.n_6_4_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_4_zpos.txt",net0.n_6_4_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_4_zneg.txt",net0.n_6_4_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_4_xpos.txt",net0.n_6_4_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_4_xneg.txt",net0.n_6_4_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_4_ypos.txt",net0.n_6_4_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_4_yneg.txt",net0.n_6_4_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_4_zpos.txt",net0.n_6_4_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_4_zneg.txt",net0.n_6_4_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_5_local.txt",net0.n_6_4_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_5_xpos.txt",net0.n_6_4_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_5_xneg.txt",net0.n_6_4_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_5_ypos.txt",net0.n_6_4_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_5_yneg.txt",net0.n_6_4_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_5_zpos.txt",net0.n_6_4_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_5_zneg.txt",net0.n_6_4_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_5_xpos.txt",net0.n_6_4_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_5_xneg.txt",net0.n_6_4_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_5_ypos.txt",net0.n_6_4_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_5_yneg.txt",net0.n_6_4_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_5_zpos.txt",net0.n_6_4_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_5_zneg.txt",net0.n_6_4_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_5_xpos.txt",net0.n_6_4_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_5_xneg.txt",net0.n_6_4_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_5_ypos.txt",net0.n_6_4_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_5_yneg.txt",net0.n_6_4_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_5_zpos.txt",net0.n_6_4_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_5_zneg.txt",net0.n_6_4_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_6_local.txt",net0.n_6_4_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_6_xpos.txt",net0.n_6_4_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_6_xneg.txt",net0.n_6_4_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_6_ypos.txt",net0.n_6_4_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_6_yneg.txt",net0.n_6_4_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_6_zpos.txt",net0.n_6_4_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_6_zneg.txt",net0.n_6_4_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_6_xpos.txt",net0.n_6_4_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_6_xneg.txt",net0.n_6_4_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_6_ypos.txt",net0.n_6_4_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_6_yneg.txt",net0.n_6_4_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_6_zpos.txt",net0.n_6_4_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_6_zneg.txt",net0.n_6_4_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_6_xpos.txt",net0.n_6_4_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_6_xneg.txt",net0.n_6_4_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_6_ypos.txt",net0.n_6_4_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_6_yneg.txt",net0.n_6_4_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_6_zpos.txt",net0.n_6_4_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_6_zneg.txt",net0.n_6_4_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_7_local.txt",net0.n_6_4_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_7_xpos.txt",net0.n_6_4_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_7_xneg.txt",net0.n_6_4_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_7_ypos.txt",net0.n_6_4_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_7_yneg.txt",net0.n_6_4_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_7_zpos.txt",net0.n_6_4_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_4_7_zneg.txt",net0.n_6_4_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_7_xpos.txt",net0.n_6_4_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_7_xneg.txt",net0.n_6_4_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_7_ypos.txt",net0.n_6_4_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_7_yneg.txt",net0.n_6_4_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_7_zpos.txt",net0.n_6_4_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_4_7_zneg.txt",net0.n_6_4_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_7_xpos.txt",net0.n_6_4_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_7_xneg.txt",net0.n_6_4_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_7_ypos.txt",net0.n_6_4_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_7_yneg.txt",net0.n_6_4_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_7_zpos.txt",net0.n_6_4_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_4_7_zneg.txt",net0.n_6_4_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_0_local.txt",net0.n_6_5_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_0_xpos.txt",net0.n_6_5_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_0_xneg.txt",net0.n_6_5_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_0_ypos.txt",net0.n_6_5_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_0_yneg.txt",net0.n_6_5_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_0_zpos.txt",net0.n_6_5_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_0_zneg.txt",net0.n_6_5_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_0_xpos.txt",net0.n_6_5_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_0_xneg.txt",net0.n_6_5_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_0_ypos.txt",net0.n_6_5_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_0_yneg.txt",net0.n_6_5_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_0_zpos.txt",net0.n_6_5_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_0_zneg.txt",net0.n_6_5_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_0_xpos.txt",net0.n_6_5_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_0_xneg.txt",net0.n_6_5_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_0_ypos.txt",net0.n_6_5_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_0_yneg.txt",net0.n_6_5_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_0_zpos.txt",net0.n_6_5_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_0_zneg.txt",net0.n_6_5_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_1_local.txt",net0.n_6_5_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_1_xpos.txt",net0.n_6_5_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_1_xneg.txt",net0.n_6_5_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_1_ypos.txt",net0.n_6_5_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_1_yneg.txt",net0.n_6_5_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_1_zpos.txt",net0.n_6_5_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_1_zneg.txt",net0.n_6_5_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_1_xpos.txt",net0.n_6_5_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_1_xneg.txt",net0.n_6_5_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_1_ypos.txt",net0.n_6_5_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_1_yneg.txt",net0.n_6_5_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_1_zpos.txt",net0.n_6_5_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_1_zneg.txt",net0.n_6_5_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_1_xpos.txt",net0.n_6_5_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_1_xneg.txt",net0.n_6_5_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_1_ypos.txt",net0.n_6_5_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_1_yneg.txt",net0.n_6_5_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_1_zpos.txt",net0.n_6_5_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_1_zneg.txt",net0.n_6_5_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_2_local.txt",net0.n_6_5_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_2_xpos.txt",net0.n_6_5_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_2_xneg.txt",net0.n_6_5_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_2_ypos.txt",net0.n_6_5_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_2_yneg.txt",net0.n_6_5_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_2_zpos.txt",net0.n_6_5_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_2_zneg.txt",net0.n_6_5_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_2_xpos.txt",net0.n_6_5_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_2_xneg.txt",net0.n_6_5_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_2_ypos.txt",net0.n_6_5_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_2_yneg.txt",net0.n_6_5_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_2_zpos.txt",net0.n_6_5_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_2_zneg.txt",net0.n_6_5_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_2_xpos.txt",net0.n_6_5_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_2_xneg.txt",net0.n_6_5_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_2_ypos.txt",net0.n_6_5_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_2_yneg.txt",net0.n_6_5_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_2_zpos.txt",net0.n_6_5_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_2_zneg.txt",net0.n_6_5_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_3_local.txt",net0.n_6_5_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_3_xpos.txt",net0.n_6_5_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_3_xneg.txt",net0.n_6_5_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_3_ypos.txt",net0.n_6_5_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_3_yneg.txt",net0.n_6_5_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_3_zpos.txt",net0.n_6_5_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_3_zneg.txt",net0.n_6_5_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_3_xpos.txt",net0.n_6_5_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_3_xneg.txt",net0.n_6_5_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_3_ypos.txt",net0.n_6_5_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_3_yneg.txt",net0.n_6_5_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_3_zpos.txt",net0.n_6_5_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_3_zneg.txt",net0.n_6_5_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_3_xpos.txt",net0.n_6_5_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_3_xneg.txt",net0.n_6_5_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_3_ypos.txt",net0.n_6_5_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_3_yneg.txt",net0.n_6_5_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_3_zpos.txt",net0.n_6_5_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_3_zneg.txt",net0.n_6_5_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_4_local.txt",net0.n_6_5_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_4_xpos.txt",net0.n_6_5_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_4_xneg.txt",net0.n_6_5_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_4_ypos.txt",net0.n_6_5_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_4_yneg.txt",net0.n_6_5_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_4_zpos.txt",net0.n_6_5_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_4_zneg.txt",net0.n_6_5_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_4_xpos.txt",net0.n_6_5_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_4_xneg.txt",net0.n_6_5_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_4_ypos.txt",net0.n_6_5_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_4_yneg.txt",net0.n_6_5_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_4_zpos.txt",net0.n_6_5_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_4_zneg.txt",net0.n_6_5_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_4_xpos.txt",net0.n_6_5_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_4_xneg.txt",net0.n_6_5_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_4_ypos.txt",net0.n_6_5_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_4_yneg.txt",net0.n_6_5_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_4_zpos.txt",net0.n_6_5_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_4_zneg.txt",net0.n_6_5_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_5_local.txt",net0.n_6_5_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_5_xpos.txt",net0.n_6_5_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_5_xneg.txt",net0.n_6_5_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_5_ypos.txt",net0.n_6_5_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_5_yneg.txt",net0.n_6_5_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_5_zpos.txt",net0.n_6_5_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_5_zneg.txt",net0.n_6_5_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_5_xpos.txt",net0.n_6_5_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_5_xneg.txt",net0.n_6_5_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_5_ypos.txt",net0.n_6_5_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_5_yneg.txt",net0.n_6_5_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_5_zpos.txt",net0.n_6_5_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_5_zneg.txt",net0.n_6_5_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_5_xpos.txt",net0.n_6_5_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_5_xneg.txt",net0.n_6_5_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_5_ypos.txt",net0.n_6_5_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_5_yneg.txt",net0.n_6_5_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_5_zpos.txt",net0.n_6_5_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_5_zneg.txt",net0.n_6_5_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_6_local.txt",net0.n_6_5_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_6_xpos.txt",net0.n_6_5_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_6_xneg.txt",net0.n_6_5_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_6_ypos.txt",net0.n_6_5_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_6_yneg.txt",net0.n_6_5_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_6_zpos.txt",net0.n_6_5_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_6_zneg.txt",net0.n_6_5_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_6_xpos.txt",net0.n_6_5_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_6_xneg.txt",net0.n_6_5_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_6_ypos.txt",net0.n_6_5_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_6_yneg.txt",net0.n_6_5_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_6_zpos.txt",net0.n_6_5_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_6_zneg.txt",net0.n_6_5_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_6_xpos.txt",net0.n_6_5_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_6_xneg.txt",net0.n_6_5_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_6_ypos.txt",net0.n_6_5_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_6_yneg.txt",net0.n_6_5_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_6_zpos.txt",net0.n_6_5_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_6_zneg.txt",net0.n_6_5_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_7_local.txt",net0.n_6_5_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_7_xpos.txt",net0.n_6_5_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_7_xneg.txt",net0.n_6_5_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_7_ypos.txt",net0.n_6_5_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_7_yneg.txt",net0.n_6_5_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_7_zpos.txt",net0.n_6_5_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_5_7_zneg.txt",net0.n_6_5_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_7_xpos.txt",net0.n_6_5_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_7_xneg.txt",net0.n_6_5_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_7_ypos.txt",net0.n_6_5_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_7_yneg.txt",net0.n_6_5_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_7_zpos.txt",net0.n_6_5_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_5_7_zneg.txt",net0.n_6_5_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_7_xpos.txt",net0.n_6_5_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_7_xneg.txt",net0.n_6_5_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_7_ypos.txt",net0.n_6_5_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_7_yneg.txt",net0.n_6_5_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_7_zpos.txt",net0.n_6_5_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_5_7_zneg.txt",net0.n_6_5_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_0_local.txt",net0.n_6_6_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_0_xpos.txt",net0.n_6_6_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_0_xneg.txt",net0.n_6_6_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_0_ypos.txt",net0.n_6_6_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_0_yneg.txt",net0.n_6_6_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_0_zpos.txt",net0.n_6_6_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_0_zneg.txt",net0.n_6_6_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_0_xpos.txt",net0.n_6_6_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_0_xneg.txt",net0.n_6_6_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_0_ypos.txt",net0.n_6_6_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_0_yneg.txt",net0.n_6_6_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_0_zpos.txt",net0.n_6_6_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_0_zneg.txt",net0.n_6_6_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_0_xpos.txt",net0.n_6_6_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_0_xneg.txt",net0.n_6_6_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_0_ypos.txt",net0.n_6_6_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_0_yneg.txt",net0.n_6_6_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_0_zpos.txt",net0.n_6_6_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_0_zneg.txt",net0.n_6_6_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_1_local.txt",net0.n_6_6_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_1_xpos.txt",net0.n_6_6_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_1_xneg.txt",net0.n_6_6_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_1_ypos.txt",net0.n_6_6_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_1_yneg.txt",net0.n_6_6_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_1_zpos.txt",net0.n_6_6_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_1_zneg.txt",net0.n_6_6_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_1_xpos.txt",net0.n_6_6_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_1_xneg.txt",net0.n_6_6_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_1_ypos.txt",net0.n_6_6_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_1_yneg.txt",net0.n_6_6_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_1_zpos.txt",net0.n_6_6_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_1_zneg.txt",net0.n_6_6_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_1_xpos.txt",net0.n_6_6_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_1_xneg.txt",net0.n_6_6_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_1_ypos.txt",net0.n_6_6_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_1_yneg.txt",net0.n_6_6_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_1_zpos.txt",net0.n_6_6_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_1_zneg.txt",net0.n_6_6_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_2_local.txt",net0.n_6_6_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_2_xpos.txt",net0.n_6_6_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_2_xneg.txt",net0.n_6_6_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_2_ypos.txt",net0.n_6_6_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_2_yneg.txt",net0.n_6_6_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_2_zpos.txt",net0.n_6_6_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_2_zneg.txt",net0.n_6_6_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_2_xpos.txt",net0.n_6_6_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_2_xneg.txt",net0.n_6_6_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_2_ypos.txt",net0.n_6_6_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_2_yneg.txt",net0.n_6_6_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_2_zpos.txt",net0.n_6_6_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_2_zneg.txt",net0.n_6_6_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_2_xpos.txt",net0.n_6_6_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_2_xneg.txt",net0.n_6_6_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_2_ypos.txt",net0.n_6_6_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_2_yneg.txt",net0.n_6_6_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_2_zpos.txt",net0.n_6_6_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_2_zneg.txt",net0.n_6_6_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_3_local.txt",net0.n_6_6_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_3_xpos.txt",net0.n_6_6_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_3_xneg.txt",net0.n_6_6_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_3_ypos.txt",net0.n_6_6_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_3_yneg.txt",net0.n_6_6_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_3_zpos.txt",net0.n_6_6_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_3_zneg.txt",net0.n_6_6_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_3_xpos.txt",net0.n_6_6_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_3_xneg.txt",net0.n_6_6_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_3_ypos.txt",net0.n_6_6_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_3_yneg.txt",net0.n_6_6_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_3_zpos.txt",net0.n_6_6_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_3_zneg.txt",net0.n_6_6_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_3_xpos.txt",net0.n_6_6_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_3_xneg.txt",net0.n_6_6_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_3_ypos.txt",net0.n_6_6_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_3_yneg.txt",net0.n_6_6_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_3_zpos.txt",net0.n_6_6_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_3_zneg.txt",net0.n_6_6_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_4_local.txt",net0.n_6_6_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_4_xpos.txt",net0.n_6_6_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_4_xneg.txt",net0.n_6_6_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_4_ypos.txt",net0.n_6_6_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_4_yneg.txt",net0.n_6_6_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_4_zpos.txt",net0.n_6_6_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_4_zneg.txt",net0.n_6_6_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_4_xpos.txt",net0.n_6_6_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_4_xneg.txt",net0.n_6_6_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_4_ypos.txt",net0.n_6_6_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_4_yneg.txt",net0.n_6_6_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_4_zpos.txt",net0.n_6_6_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_4_zneg.txt",net0.n_6_6_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_4_xpos.txt",net0.n_6_6_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_4_xneg.txt",net0.n_6_6_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_4_ypos.txt",net0.n_6_6_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_4_yneg.txt",net0.n_6_6_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_4_zpos.txt",net0.n_6_6_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_4_zneg.txt",net0.n_6_6_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_5_local.txt",net0.n_6_6_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_5_xpos.txt",net0.n_6_6_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_5_xneg.txt",net0.n_6_6_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_5_ypos.txt",net0.n_6_6_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_5_yneg.txt",net0.n_6_6_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_5_zpos.txt",net0.n_6_6_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_5_zneg.txt",net0.n_6_6_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_5_xpos.txt",net0.n_6_6_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_5_xneg.txt",net0.n_6_6_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_5_ypos.txt",net0.n_6_6_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_5_yneg.txt",net0.n_6_6_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_5_zpos.txt",net0.n_6_6_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_5_zneg.txt",net0.n_6_6_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_5_xpos.txt",net0.n_6_6_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_5_xneg.txt",net0.n_6_6_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_5_ypos.txt",net0.n_6_6_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_5_yneg.txt",net0.n_6_6_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_5_zpos.txt",net0.n_6_6_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_5_zneg.txt",net0.n_6_6_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_6_local.txt",net0.n_6_6_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_6_xpos.txt",net0.n_6_6_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_6_xneg.txt",net0.n_6_6_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_6_ypos.txt",net0.n_6_6_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_6_yneg.txt",net0.n_6_6_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_6_zpos.txt",net0.n_6_6_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_6_zneg.txt",net0.n_6_6_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_6_xpos.txt",net0.n_6_6_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_6_xneg.txt",net0.n_6_6_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_6_ypos.txt",net0.n_6_6_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_6_yneg.txt",net0.n_6_6_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_6_zpos.txt",net0.n_6_6_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_6_zneg.txt",net0.n_6_6_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_6_xpos.txt",net0.n_6_6_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_6_xneg.txt",net0.n_6_6_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_6_ypos.txt",net0.n_6_6_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_6_yneg.txt",net0.n_6_6_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_6_zpos.txt",net0.n_6_6_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_6_zneg.txt",net0.n_6_6_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_7_local.txt",net0.n_6_6_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_7_xpos.txt",net0.n_6_6_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_7_xneg.txt",net0.n_6_6_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_7_ypos.txt",net0.n_6_6_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_7_yneg.txt",net0.n_6_6_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_7_zpos.txt",net0.n_6_6_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_6_7_zneg.txt",net0.n_6_6_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_7_xpos.txt",net0.n_6_6_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_7_xneg.txt",net0.n_6_6_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_7_ypos.txt",net0.n_6_6_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_7_yneg.txt",net0.n_6_6_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_7_zpos.txt",net0.n_6_6_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_6_7_zneg.txt",net0.n_6_6_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_7_xpos.txt",net0.n_6_6_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_7_xneg.txt",net0.n_6_6_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_7_ypos.txt",net0.n_6_6_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_7_yneg.txt",net0.n_6_6_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_7_zpos.txt",net0.n_6_6_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_6_7_zneg.txt",net0.n_6_6_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_0_local.txt",net0.n_6_7_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_0_xpos.txt",net0.n_6_7_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_0_xneg.txt",net0.n_6_7_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_0_ypos.txt",net0.n_6_7_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_0_yneg.txt",net0.n_6_7_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_0_zpos.txt",net0.n_6_7_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_0_zneg.txt",net0.n_6_7_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_0_xpos.txt",net0.n_6_7_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_0_xneg.txt",net0.n_6_7_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_0_ypos.txt",net0.n_6_7_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_0_yneg.txt",net0.n_6_7_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_0_zpos.txt",net0.n_6_7_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_0_zneg.txt",net0.n_6_7_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_0_xpos.txt",net0.n_6_7_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_0_xneg.txt",net0.n_6_7_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_0_ypos.txt",net0.n_6_7_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_0_yneg.txt",net0.n_6_7_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_0_zpos.txt",net0.n_6_7_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_0_zneg.txt",net0.n_6_7_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_1_local.txt",net0.n_6_7_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_1_xpos.txt",net0.n_6_7_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_1_xneg.txt",net0.n_6_7_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_1_ypos.txt",net0.n_6_7_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_1_yneg.txt",net0.n_6_7_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_1_zpos.txt",net0.n_6_7_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_1_zneg.txt",net0.n_6_7_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_1_xpos.txt",net0.n_6_7_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_1_xneg.txt",net0.n_6_7_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_1_ypos.txt",net0.n_6_7_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_1_yneg.txt",net0.n_6_7_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_1_zpos.txt",net0.n_6_7_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_1_zneg.txt",net0.n_6_7_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_1_xpos.txt",net0.n_6_7_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_1_xneg.txt",net0.n_6_7_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_1_ypos.txt",net0.n_6_7_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_1_yneg.txt",net0.n_6_7_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_1_zpos.txt",net0.n_6_7_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_1_zneg.txt",net0.n_6_7_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_2_local.txt",net0.n_6_7_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_2_xpos.txt",net0.n_6_7_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_2_xneg.txt",net0.n_6_7_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_2_ypos.txt",net0.n_6_7_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_2_yneg.txt",net0.n_6_7_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_2_zpos.txt",net0.n_6_7_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_2_zneg.txt",net0.n_6_7_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_2_xpos.txt",net0.n_6_7_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_2_xneg.txt",net0.n_6_7_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_2_ypos.txt",net0.n_6_7_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_2_yneg.txt",net0.n_6_7_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_2_zpos.txt",net0.n_6_7_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_2_zneg.txt",net0.n_6_7_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_2_xpos.txt",net0.n_6_7_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_2_xneg.txt",net0.n_6_7_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_2_ypos.txt",net0.n_6_7_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_2_yneg.txt",net0.n_6_7_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_2_zpos.txt",net0.n_6_7_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_2_zneg.txt",net0.n_6_7_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_3_local.txt",net0.n_6_7_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_3_xpos.txt",net0.n_6_7_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_3_xneg.txt",net0.n_6_7_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_3_ypos.txt",net0.n_6_7_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_3_yneg.txt",net0.n_6_7_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_3_zpos.txt",net0.n_6_7_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_3_zneg.txt",net0.n_6_7_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_3_xpos.txt",net0.n_6_7_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_3_xneg.txt",net0.n_6_7_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_3_ypos.txt",net0.n_6_7_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_3_yneg.txt",net0.n_6_7_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_3_zpos.txt",net0.n_6_7_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_3_zneg.txt",net0.n_6_7_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_3_xpos.txt",net0.n_6_7_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_3_xneg.txt",net0.n_6_7_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_3_ypos.txt",net0.n_6_7_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_3_yneg.txt",net0.n_6_7_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_3_zpos.txt",net0.n_6_7_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_3_zneg.txt",net0.n_6_7_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_4_local.txt",net0.n_6_7_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_4_xpos.txt",net0.n_6_7_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_4_xneg.txt",net0.n_6_7_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_4_ypos.txt",net0.n_6_7_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_4_yneg.txt",net0.n_6_7_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_4_zpos.txt",net0.n_6_7_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_4_zneg.txt",net0.n_6_7_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_4_xpos.txt",net0.n_6_7_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_4_xneg.txt",net0.n_6_7_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_4_ypos.txt",net0.n_6_7_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_4_yneg.txt",net0.n_6_7_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_4_zpos.txt",net0.n_6_7_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_4_zneg.txt",net0.n_6_7_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_4_xpos.txt",net0.n_6_7_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_4_xneg.txt",net0.n_6_7_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_4_ypos.txt",net0.n_6_7_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_4_yneg.txt",net0.n_6_7_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_4_zpos.txt",net0.n_6_7_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_4_zneg.txt",net0.n_6_7_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_5_local.txt",net0.n_6_7_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_5_xpos.txt",net0.n_6_7_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_5_xneg.txt",net0.n_6_7_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_5_ypos.txt",net0.n_6_7_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_5_yneg.txt",net0.n_6_7_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_5_zpos.txt",net0.n_6_7_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_5_zneg.txt",net0.n_6_7_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_5_xpos.txt",net0.n_6_7_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_5_xneg.txt",net0.n_6_7_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_5_ypos.txt",net0.n_6_7_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_5_yneg.txt",net0.n_6_7_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_5_zpos.txt",net0.n_6_7_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_5_zneg.txt",net0.n_6_7_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_5_xpos.txt",net0.n_6_7_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_5_xneg.txt",net0.n_6_7_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_5_ypos.txt",net0.n_6_7_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_5_yneg.txt",net0.n_6_7_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_5_zpos.txt",net0.n_6_7_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_5_zneg.txt",net0.n_6_7_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_6_local.txt",net0.n_6_7_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_6_xpos.txt",net0.n_6_7_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_6_xneg.txt",net0.n_6_7_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_6_ypos.txt",net0.n_6_7_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_6_yneg.txt",net0.n_6_7_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_6_zpos.txt",net0.n_6_7_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_6_zneg.txt",net0.n_6_7_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_6_xpos.txt",net0.n_6_7_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_6_xneg.txt",net0.n_6_7_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_6_ypos.txt",net0.n_6_7_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_6_yneg.txt",net0.n_6_7_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_6_zpos.txt",net0.n_6_7_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_6_zneg.txt",net0.n_6_7_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_6_xpos.txt",net0.n_6_7_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_6_xneg.txt",net0.n_6_7_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_6_ypos.txt",net0.n_6_7_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_6_yneg.txt",net0.n_6_7_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_6_zpos.txt",net0.n_6_7_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_6_zneg.txt",net0.n_6_7_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_7_local.txt",net0.n_6_7_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_7_xpos.txt",net0.n_6_7_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_7_xneg.txt",net0.n_6_7_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_7_ypos.txt",net0.n_6_7_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_7_yneg.txt",net0.n_6_7_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_7_zpos.txt",net0.n_6_7_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_6_7_7_zneg.txt",net0.n_6_7_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_7_xpos.txt",net0.n_6_7_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_7_xneg.txt",net0.n_6_7_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_7_ypos.txt",net0.n_6_7_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_7_yneg.txt",net0.n_6_7_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_7_zpos.txt",net0.n_6_7_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_6_7_7_zneg.txt",net0.n_6_7_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_7_xpos.txt",net0.n_6_7_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_7_xneg.txt",net0.n_6_7_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_7_ypos.txt",net0.n_6_7_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_7_yneg.txt",net0.n_6_7_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_7_zpos.txt",net0.n_6_7_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_6_7_7_zneg.txt",net0.n_6_7_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_0_local.txt",net0.n_7_0_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_0_xpos.txt",net0.n_7_0_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_0_xneg.txt",net0.n_7_0_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_0_ypos.txt",net0.n_7_0_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_0_yneg.txt",net0.n_7_0_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_0_zpos.txt",net0.n_7_0_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_0_zneg.txt",net0.n_7_0_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_0_xpos.txt",net0.n_7_0_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_0_xneg.txt",net0.n_7_0_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_0_ypos.txt",net0.n_7_0_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_0_yneg.txt",net0.n_7_0_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_0_zpos.txt",net0.n_7_0_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_0_zneg.txt",net0.n_7_0_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_0_xpos.txt",net0.n_7_0_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_0_xneg.txt",net0.n_7_0_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_0_ypos.txt",net0.n_7_0_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_0_yneg.txt",net0.n_7_0_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_0_zpos.txt",net0.n_7_0_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_0_zneg.txt",net0.n_7_0_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_1_local.txt",net0.n_7_0_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_1_xpos.txt",net0.n_7_0_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_1_xneg.txt",net0.n_7_0_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_1_ypos.txt",net0.n_7_0_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_1_yneg.txt",net0.n_7_0_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_1_zpos.txt",net0.n_7_0_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_1_zneg.txt",net0.n_7_0_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_1_xpos.txt",net0.n_7_0_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_1_xneg.txt",net0.n_7_0_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_1_ypos.txt",net0.n_7_0_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_1_yneg.txt",net0.n_7_0_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_1_zpos.txt",net0.n_7_0_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_1_zneg.txt",net0.n_7_0_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_1_xpos.txt",net0.n_7_0_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_1_xneg.txt",net0.n_7_0_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_1_ypos.txt",net0.n_7_0_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_1_yneg.txt",net0.n_7_0_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_1_zpos.txt",net0.n_7_0_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_1_zneg.txt",net0.n_7_0_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_2_local.txt",net0.n_7_0_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_2_xpos.txt",net0.n_7_0_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_2_xneg.txt",net0.n_7_0_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_2_ypos.txt",net0.n_7_0_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_2_yneg.txt",net0.n_7_0_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_2_zpos.txt",net0.n_7_0_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_2_zneg.txt",net0.n_7_0_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_2_xpos.txt",net0.n_7_0_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_2_xneg.txt",net0.n_7_0_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_2_ypos.txt",net0.n_7_0_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_2_yneg.txt",net0.n_7_0_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_2_zpos.txt",net0.n_7_0_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_2_zneg.txt",net0.n_7_0_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_2_xpos.txt",net0.n_7_0_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_2_xneg.txt",net0.n_7_0_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_2_ypos.txt",net0.n_7_0_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_2_yneg.txt",net0.n_7_0_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_2_zpos.txt",net0.n_7_0_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_2_zneg.txt",net0.n_7_0_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_3_local.txt",net0.n_7_0_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_3_xpos.txt",net0.n_7_0_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_3_xneg.txt",net0.n_7_0_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_3_ypos.txt",net0.n_7_0_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_3_yneg.txt",net0.n_7_0_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_3_zpos.txt",net0.n_7_0_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_3_zneg.txt",net0.n_7_0_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_3_xpos.txt",net0.n_7_0_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_3_xneg.txt",net0.n_7_0_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_3_ypos.txt",net0.n_7_0_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_3_yneg.txt",net0.n_7_0_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_3_zpos.txt",net0.n_7_0_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_3_zneg.txt",net0.n_7_0_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_3_xpos.txt",net0.n_7_0_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_3_xneg.txt",net0.n_7_0_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_3_ypos.txt",net0.n_7_0_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_3_yneg.txt",net0.n_7_0_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_3_zpos.txt",net0.n_7_0_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_3_zneg.txt",net0.n_7_0_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_4_local.txt",net0.n_7_0_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_4_xpos.txt",net0.n_7_0_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_4_xneg.txt",net0.n_7_0_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_4_ypos.txt",net0.n_7_0_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_4_yneg.txt",net0.n_7_0_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_4_zpos.txt",net0.n_7_0_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_4_zneg.txt",net0.n_7_0_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_4_xpos.txt",net0.n_7_0_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_4_xneg.txt",net0.n_7_0_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_4_ypos.txt",net0.n_7_0_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_4_yneg.txt",net0.n_7_0_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_4_zpos.txt",net0.n_7_0_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_4_zneg.txt",net0.n_7_0_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_4_xpos.txt",net0.n_7_0_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_4_xneg.txt",net0.n_7_0_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_4_ypos.txt",net0.n_7_0_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_4_yneg.txt",net0.n_7_0_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_4_zpos.txt",net0.n_7_0_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_4_zneg.txt",net0.n_7_0_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_5_local.txt",net0.n_7_0_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_5_xpos.txt",net0.n_7_0_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_5_xneg.txt",net0.n_7_0_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_5_ypos.txt",net0.n_7_0_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_5_yneg.txt",net0.n_7_0_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_5_zpos.txt",net0.n_7_0_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_5_zneg.txt",net0.n_7_0_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_5_xpos.txt",net0.n_7_0_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_5_xneg.txt",net0.n_7_0_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_5_ypos.txt",net0.n_7_0_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_5_yneg.txt",net0.n_7_0_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_5_zpos.txt",net0.n_7_0_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_5_zneg.txt",net0.n_7_0_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_5_xpos.txt",net0.n_7_0_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_5_xneg.txt",net0.n_7_0_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_5_ypos.txt",net0.n_7_0_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_5_yneg.txt",net0.n_7_0_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_5_zpos.txt",net0.n_7_0_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_5_zneg.txt",net0.n_7_0_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_6_local.txt",net0.n_7_0_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_6_xpos.txt",net0.n_7_0_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_6_xneg.txt",net0.n_7_0_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_6_ypos.txt",net0.n_7_0_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_6_yneg.txt",net0.n_7_0_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_6_zpos.txt",net0.n_7_0_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_6_zneg.txt",net0.n_7_0_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_6_xpos.txt",net0.n_7_0_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_6_xneg.txt",net0.n_7_0_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_6_ypos.txt",net0.n_7_0_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_6_yneg.txt",net0.n_7_0_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_6_zpos.txt",net0.n_7_0_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_6_zneg.txt",net0.n_7_0_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_6_xpos.txt",net0.n_7_0_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_6_xneg.txt",net0.n_7_0_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_6_ypos.txt",net0.n_7_0_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_6_yneg.txt",net0.n_7_0_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_6_zpos.txt",net0.n_7_0_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_6_zneg.txt",net0.n_7_0_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_7_local.txt",net0.n_7_0_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_7_xpos.txt",net0.n_7_0_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_7_xneg.txt",net0.n_7_0_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_7_ypos.txt",net0.n_7_0_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_7_yneg.txt",net0.n_7_0_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_7_zpos.txt",net0.n_7_0_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_0_7_zneg.txt",net0.n_7_0_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_7_xpos.txt",net0.n_7_0_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_7_xneg.txt",net0.n_7_0_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_7_ypos.txt",net0.n_7_0_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_7_yneg.txt",net0.n_7_0_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_7_zpos.txt",net0.n_7_0_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_0_7_zneg.txt",net0.n_7_0_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_7_xpos.txt",net0.n_7_0_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_7_xneg.txt",net0.n_7_0_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_7_ypos.txt",net0.n_7_0_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_7_yneg.txt",net0.n_7_0_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_7_zpos.txt",net0.n_7_0_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_0_7_zneg.txt",net0.n_7_0_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_0_local.txt",net0.n_7_1_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_0_xpos.txt",net0.n_7_1_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_0_xneg.txt",net0.n_7_1_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_0_ypos.txt",net0.n_7_1_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_0_yneg.txt",net0.n_7_1_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_0_zpos.txt",net0.n_7_1_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_0_zneg.txt",net0.n_7_1_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_0_xpos.txt",net0.n_7_1_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_0_xneg.txt",net0.n_7_1_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_0_ypos.txt",net0.n_7_1_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_0_yneg.txt",net0.n_7_1_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_0_zpos.txt",net0.n_7_1_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_0_zneg.txt",net0.n_7_1_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_0_xpos.txt",net0.n_7_1_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_0_xneg.txt",net0.n_7_1_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_0_ypos.txt",net0.n_7_1_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_0_yneg.txt",net0.n_7_1_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_0_zpos.txt",net0.n_7_1_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_0_zneg.txt",net0.n_7_1_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_1_local.txt",net0.n_7_1_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_1_xpos.txt",net0.n_7_1_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_1_xneg.txt",net0.n_7_1_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_1_ypos.txt",net0.n_7_1_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_1_yneg.txt",net0.n_7_1_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_1_zpos.txt",net0.n_7_1_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_1_zneg.txt",net0.n_7_1_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_1_xpos.txt",net0.n_7_1_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_1_xneg.txt",net0.n_7_1_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_1_ypos.txt",net0.n_7_1_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_1_yneg.txt",net0.n_7_1_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_1_zpos.txt",net0.n_7_1_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_1_zneg.txt",net0.n_7_1_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_1_xpos.txt",net0.n_7_1_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_1_xneg.txt",net0.n_7_1_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_1_ypos.txt",net0.n_7_1_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_1_yneg.txt",net0.n_7_1_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_1_zpos.txt",net0.n_7_1_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_1_zneg.txt",net0.n_7_1_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_2_local.txt",net0.n_7_1_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_2_xpos.txt",net0.n_7_1_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_2_xneg.txt",net0.n_7_1_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_2_ypos.txt",net0.n_7_1_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_2_yneg.txt",net0.n_7_1_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_2_zpos.txt",net0.n_7_1_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_2_zneg.txt",net0.n_7_1_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_2_xpos.txt",net0.n_7_1_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_2_xneg.txt",net0.n_7_1_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_2_ypos.txt",net0.n_7_1_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_2_yneg.txt",net0.n_7_1_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_2_zpos.txt",net0.n_7_1_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_2_zneg.txt",net0.n_7_1_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_2_xpos.txt",net0.n_7_1_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_2_xneg.txt",net0.n_7_1_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_2_ypos.txt",net0.n_7_1_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_2_yneg.txt",net0.n_7_1_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_2_zpos.txt",net0.n_7_1_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_2_zneg.txt",net0.n_7_1_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_3_local.txt",net0.n_7_1_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_3_xpos.txt",net0.n_7_1_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_3_xneg.txt",net0.n_7_1_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_3_ypos.txt",net0.n_7_1_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_3_yneg.txt",net0.n_7_1_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_3_zpos.txt",net0.n_7_1_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_3_zneg.txt",net0.n_7_1_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_3_xpos.txt",net0.n_7_1_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_3_xneg.txt",net0.n_7_1_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_3_ypos.txt",net0.n_7_1_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_3_yneg.txt",net0.n_7_1_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_3_zpos.txt",net0.n_7_1_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_3_zneg.txt",net0.n_7_1_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_3_xpos.txt",net0.n_7_1_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_3_xneg.txt",net0.n_7_1_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_3_ypos.txt",net0.n_7_1_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_3_yneg.txt",net0.n_7_1_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_3_zpos.txt",net0.n_7_1_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_3_zneg.txt",net0.n_7_1_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_4_local.txt",net0.n_7_1_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_4_xpos.txt",net0.n_7_1_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_4_xneg.txt",net0.n_7_1_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_4_ypos.txt",net0.n_7_1_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_4_yneg.txt",net0.n_7_1_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_4_zpos.txt",net0.n_7_1_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_4_zneg.txt",net0.n_7_1_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_4_xpos.txt",net0.n_7_1_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_4_xneg.txt",net0.n_7_1_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_4_ypos.txt",net0.n_7_1_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_4_yneg.txt",net0.n_7_1_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_4_zpos.txt",net0.n_7_1_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_4_zneg.txt",net0.n_7_1_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_4_xpos.txt",net0.n_7_1_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_4_xneg.txt",net0.n_7_1_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_4_ypos.txt",net0.n_7_1_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_4_yneg.txt",net0.n_7_1_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_4_zpos.txt",net0.n_7_1_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_4_zneg.txt",net0.n_7_1_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_5_local.txt",net0.n_7_1_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_5_xpos.txt",net0.n_7_1_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_5_xneg.txt",net0.n_7_1_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_5_ypos.txt",net0.n_7_1_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_5_yneg.txt",net0.n_7_1_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_5_zpos.txt",net0.n_7_1_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_5_zneg.txt",net0.n_7_1_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_5_xpos.txt",net0.n_7_1_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_5_xneg.txt",net0.n_7_1_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_5_ypos.txt",net0.n_7_1_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_5_yneg.txt",net0.n_7_1_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_5_zpos.txt",net0.n_7_1_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_5_zneg.txt",net0.n_7_1_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_5_xpos.txt",net0.n_7_1_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_5_xneg.txt",net0.n_7_1_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_5_ypos.txt",net0.n_7_1_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_5_yneg.txt",net0.n_7_1_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_5_zpos.txt",net0.n_7_1_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_5_zneg.txt",net0.n_7_1_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_6_local.txt",net0.n_7_1_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_6_xpos.txt",net0.n_7_1_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_6_xneg.txt",net0.n_7_1_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_6_ypos.txt",net0.n_7_1_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_6_yneg.txt",net0.n_7_1_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_6_zpos.txt",net0.n_7_1_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_6_zneg.txt",net0.n_7_1_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_6_xpos.txt",net0.n_7_1_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_6_xneg.txt",net0.n_7_1_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_6_ypos.txt",net0.n_7_1_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_6_yneg.txt",net0.n_7_1_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_6_zpos.txt",net0.n_7_1_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_6_zneg.txt",net0.n_7_1_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_6_xpos.txt",net0.n_7_1_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_6_xneg.txt",net0.n_7_1_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_6_ypos.txt",net0.n_7_1_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_6_yneg.txt",net0.n_7_1_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_6_zpos.txt",net0.n_7_1_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_6_zneg.txt",net0.n_7_1_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_7_local.txt",net0.n_7_1_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_7_xpos.txt",net0.n_7_1_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_7_xneg.txt",net0.n_7_1_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_7_ypos.txt",net0.n_7_1_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_7_yneg.txt",net0.n_7_1_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_7_zpos.txt",net0.n_7_1_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_1_7_zneg.txt",net0.n_7_1_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_7_xpos.txt",net0.n_7_1_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_7_xneg.txt",net0.n_7_1_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_7_ypos.txt",net0.n_7_1_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_7_yneg.txt",net0.n_7_1_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_7_zpos.txt",net0.n_7_1_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_1_7_zneg.txt",net0.n_7_1_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_7_xpos.txt",net0.n_7_1_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_7_xneg.txt",net0.n_7_1_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_7_ypos.txt",net0.n_7_1_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_7_yneg.txt",net0.n_7_1_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_7_zpos.txt",net0.n_7_1_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_1_7_zneg.txt",net0.n_7_1_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_0_local.txt",net0.n_7_2_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_0_xpos.txt",net0.n_7_2_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_0_xneg.txt",net0.n_7_2_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_0_ypos.txt",net0.n_7_2_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_0_yneg.txt",net0.n_7_2_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_0_zpos.txt",net0.n_7_2_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_0_zneg.txt",net0.n_7_2_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_0_xpos.txt",net0.n_7_2_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_0_xneg.txt",net0.n_7_2_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_0_ypos.txt",net0.n_7_2_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_0_yneg.txt",net0.n_7_2_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_0_zpos.txt",net0.n_7_2_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_0_zneg.txt",net0.n_7_2_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_0_xpos.txt",net0.n_7_2_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_0_xneg.txt",net0.n_7_2_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_0_ypos.txt",net0.n_7_2_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_0_yneg.txt",net0.n_7_2_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_0_zpos.txt",net0.n_7_2_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_0_zneg.txt",net0.n_7_2_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_1_local.txt",net0.n_7_2_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_1_xpos.txt",net0.n_7_2_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_1_xneg.txt",net0.n_7_2_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_1_ypos.txt",net0.n_7_2_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_1_yneg.txt",net0.n_7_2_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_1_zpos.txt",net0.n_7_2_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_1_zneg.txt",net0.n_7_2_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_1_xpos.txt",net0.n_7_2_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_1_xneg.txt",net0.n_7_2_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_1_ypos.txt",net0.n_7_2_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_1_yneg.txt",net0.n_7_2_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_1_zpos.txt",net0.n_7_2_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_1_zneg.txt",net0.n_7_2_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_1_xpos.txt",net0.n_7_2_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_1_xneg.txt",net0.n_7_2_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_1_ypos.txt",net0.n_7_2_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_1_yneg.txt",net0.n_7_2_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_1_zpos.txt",net0.n_7_2_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_1_zneg.txt",net0.n_7_2_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_2_local.txt",net0.n_7_2_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_2_xpos.txt",net0.n_7_2_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_2_xneg.txt",net0.n_7_2_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_2_ypos.txt",net0.n_7_2_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_2_yneg.txt",net0.n_7_2_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_2_zpos.txt",net0.n_7_2_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_2_zneg.txt",net0.n_7_2_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_2_xpos.txt",net0.n_7_2_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_2_xneg.txt",net0.n_7_2_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_2_ypos.txt",net0.n_7_2_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_2_yneg.txt",net0.n_7_2_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_2_zpos.txt",net0.n_7_2_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_2_zneg.txt",net0.n_7_2_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_2_xpos.txt",net0.n_7_2_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_2_xneg.txt",net0.n_7_2_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_2_ypos.txt",net0.n_7_2_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_2_yneg.txt",net0.n_7_2_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_2_zpos.txt",net0.n_7_2_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_2_zneg.txt",net0.n_7_2_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_3_local.txt",net0.n_7_2_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_3_xpos.txt",net0.n_7_2_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_3_xneg.txt",net0.n_7_2_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_3_ypos.txt",net0.n_7_2_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_3_yneg.txt",net0.n_7_2_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_3_zpos.txt",net0.n_7_2_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_3_zneg.txt",net0.n_7_2_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_3_xpos.txt",net0.n_7_2_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_3_xneg.txt",net0.n_7_2_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_3_ypos.txt",net0.n_7_2_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_3_yneg.txt",net0.n_7_2_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_3_zpos.txt",net0.n_7_2_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_3_zneg.txt",net0.n_7_2_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_3_xpos.txt",net0.n_7_2_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_3_xneg.txt",net0.n_7_2_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_3_ypos.txt",net0.n_7_2_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_3_yneg.txt",net0.n_7_2_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_3_zpos.txt",net0.n_7_2_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_3_zneg.txt",net0.n_7_2_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_4_local.txt",net0.n_7_2_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_4_xpos.txt",net0.n_7_2_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_4_xneg.txt",net0.n_7_2_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_4_ypos.txt",net0.n_7_2_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_4_yneg.txt",net0.n_7_2_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_4_zpos.txt",net0.n_7_2_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_4_zneg.txt",net0.n_7_2_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_4_xpos.txt",net0.n_7_2_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_4_xneg.txt",net0.n_7_2_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_4_ypos.txt",net0.n_7_2_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_4_yneg.txt",net0.n_7_2_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_4_zpos.txt",net0.n_7_2_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_4_zneg.txt",net0.n_7_2_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_4_xpos.txt",net0.n_7_2_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_4_xneg.txt",net0.n_7_2_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_4_ypos.txt",net0.n_7_2_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_4_yneg.txt",net0.n_7_2_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_4_zpos.txt",net0.n_7_2_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_4_zneg.txt",net0.n_7_2_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_5_local.txt",net0.n_7_2_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_5_xpos.txt",net0.n_7_2_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_5_xneg.txt",net0.n_7_2_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_5_ypos.txt",net0.n_7_2_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_5_yneg.txt",net0.n_7_2_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_5_zpos.txt",net0.n_7_2_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_5_zneg.txt",net0.n_7_2_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_5_xpos.txt",net0.n_7_2_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_5_xneg.txt",net0.n_7_2_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_5_ypos.txt",net0.n_7_2_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_5_yneg.txt",net0.n_7_2_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_5_zpos.txt",net0.n_7_2_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_5_zneg.txt",net0.n_7_2_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_5_xpos.txt",net0.n_7_2_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_5_xneg.txt",net0.n_7_2_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_5_ypos.txt",net0.n_7_2_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_5_yneg.txt",net0.n_7_2_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_5_zpos.txt",net0.n_7_2_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_5_zneg.txt",net0.n_7_2_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_6_local.txt",net0.n_7_2_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_6_xpos.txt",net0.n_7_2_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_6_xneg.txt",net0.n_7_2_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_6_ypos.txt",net0.n_7_2_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_6_yneg.txt",net0.n_7_2_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_6_zpos.txt",net0.n_7_2_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_6_zneg.txt",net0.n_7_2_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_6_xpos.txt",net0.n_7_2_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_6_xneg.txt",net0.n_7_2_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_6_ypos.txt",net0.n_7_2_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_6_yneg.txt",net0.n_7_2_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_6_zpos.txt",net0.n_7_2_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_6_zneg.txt",net0.n_7_2_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_6_xpos.txt",net0.n_7_2_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_6_xneg.txt",net0.n_7_2_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_6_ypos.txt",net0.n_7_2_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_6_yneg.txt",net0.n_7_2_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_6_zpos.txt",net0.n_7_2_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_6_zneg.txt",net0.n_7_2_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_7_local.txt",net0.n_7_2_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_7_xpos.txt",net0.n_7_2_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_7_xneg.txt",net0.n_7_2_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_7_ypos.txt",net0.n_7_2_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_7_yneg.txt",net0.n_7_2_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_7_zpos.txt",net0.n_7_2_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_2_7_zneg.txt",net0.n_7_2_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_7_xpos.txt",net0.n_7_2_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_7_xneg.txt",net0.n_7_2_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_7_ypos.txt",net0.n_7_2_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_7_yneg.txt",net0.n_7_2_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_7_zpos.txt",net0.n_7_2_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_2_7_zneg.txt",net0.n_7_2_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_7_xpos.txt",net0.n_7_2_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_7_xneg.txt",net0.n_7_2_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_7_ypos.txt",net0.n_7_2_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_7_yneg.txt",net0.n_7_2_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_7_zpos.txt",net0.n_7_2_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_2_7_zneg.txt",net0.n_7_2_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_0_local.txt",net0.n_7_3_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_0_xpos.txt",net0.n_7_3_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_0_xneg.txt",net0.n_7_3_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_0_ypos.txt",net0.n_7_3_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_0_yneg.txt",net0.n_7_3_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_0_zpos.txt",net0.n_7_3_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_0_zneg.txt",net0.n_7_3_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_0_xpos.txt",net0.n_7_3_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_0_xneg.txt",net0.n_7_3_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_0_ypos.txt",net0.n_7_3_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_0_yneg.txt",net0.n_7_3_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_0_zpos.txt",net0.n_7_3_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_0_zneg.txt",net0.n_7_3_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_0_xpos.txt",net0.n_7_3_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_0_xneg.txt",net0.n_7_3_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_0_ypos.txt",net0.n_7_3_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_0_yneg.txt",net0.n_7_3_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_0_zpos.txt",net0.n_7_3_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_0_zneg.txt",net0.n_7_3_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_1_local.txt",net0.n_7_3_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_1_xpos.txt",net0.n_7_3_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_1_xneg.txt",net0.n_7_3_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_1_ypos.txt",net0.n_7_3_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_1_yneg.txt",net0.n_7_3_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_1_zpos.txt",net0.n_7_3_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_1_zneg.txt",net0.n_7_3_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_1_xpos.txt",net0.n_7_3_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_1_xneg.txt",net0.n_7_3_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_1_ypos.txt",net0.n_7_3_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_1_yneg.txt",net0.n_7_3_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_1_zpos.txt",net0.n_7_3_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_1_zneg.txt",net0.n_7_3_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_1_xpos.txt",net0.n_7_3_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_1_xneg.txt",net0.n_7_3_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_1_ypos.txt",net0.n_7_3_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_1_yneg.txt",net0.n_7_3_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_1_zpos.txt",net0.n_7_3_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_1_zneg.txt",net0.n_7_3_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_2_local.txt",net0.n_7_3_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_2_xpos.txt",net0.n_7_3_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_2_xneg.txt",net0.n_7_3_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_2_ypos.txt",net0.n_7_3_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_2_yneg.txt",net0.n_7_3_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_2_zpos.txt",net0.n_7_3_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_2_zneg.txt",net0.n_7_3_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_2_xpos.txt",net0.n_7_3_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_2_xneg.txt",net0.n_7_3_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_2_ypos.txt",net0.n_7_3_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_2_yneg.txt",net0.n_7_3_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_2_zpos.txt",net0.n_7_3_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_2_zneg.txt",net0.n_7_3_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_2_xpos.txt",net0.n_7_3_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_2_xneg.txt",net0.n_7_3_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_2_ypos.txt",net0.n_7_3_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_2_yneg.txt",net0.n_7_3_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_2_zpos.txt",net0.n_7_3_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_2_zneg.txt",net0.n_7_3_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_3_local.txt",net0.n_7_3_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_3_xpos.txt",net0.n_7_3_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_3_xneg.txt",net0.n_7_3_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_3_ypos.txt",net0.n_7_3_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_3_yneg.txt",net0.n_7_3_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_3_zpos.txt",net0.n_7_3_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_3_zneg.txt",net0.n_7_3_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_3_xpos.txt",net0.n_7_3_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_3_xneg.txt",net0.n_7_3_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_3_ypos.txt",net0.n_7_3_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_3_yneg.txt",net0.n_7_3_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_3_zpos.txt",net0.n_7_3_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_3_zneg.txt",net0.n_7_3_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_3_xpos.txt",net0.n_7_3_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_3_xneg.txt",net0.n_7_3_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_3_ypos.txt",net0.n_7_3_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_3_yneg.txt",net0.n_7_3_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_3_zpos.txt",net0.n_7_3_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_3_zneg.txt",net0.n_7_3_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_4_local.txt",net0.n_7_3_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_4_xpos.txt",net0.n_7_3_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_4_xneg.txt",net0.n_7_3_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_4_ypos.txt",net0.n_7_3_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_4_yneg.txt",net0.n_7_3_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_4_zpos.txt",net0.n_7_3_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_4_zneg.txt",net0.n_7_3_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_4_xpos.txt",net0.n_7_3_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_4_xneg.txt",net0.n_7_3_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_4_ypos.txt",net0.n_7_3_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_4_yneg.txt",net0.n_7_3_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_4_zpos.txt",net0.n_7_3_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_4_zneg.txt",net0.n_7_3_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_4_xpos.txt",net0.n_7_3_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_4_xneg.txt",net0.n_7_3_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_4_ypos.txt",net0.n_7_3_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_4_yneg.txt",net0.n_7_3_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_4_zpos.txt",net0.n_7_3_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_4_zneg.txt",net0.n_7_3_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_5_local.txt",net0.n_7_3_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_5_xpos.txt",net0.n_7_3_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_5_xneg.txt",net0.n_7_3_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_5_ypos.txt",net0.n_7_3_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_5_yneg.txt",net0.n_7_3_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_5_zpos.txt",net0.n_7_3_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_5_zneg.txt",net0.n_7_3_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_5_xpos.txt",net0.n_7_3_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_5_xneg.txt",net0.n_7_3_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_5_ypos.txt",net0.n_7_3_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_5_yneg.txt",net0.n_7_3_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_5_zpos.txt",net0.n_7_3_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_5_zneg.txt",net0.n_7_3_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_5_xpos.txt",net0.n_7_3_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_5_xneg.txt",net0.n_7_3_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_5_ypos.txt",net0.n_7_3_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_5_yneg.txt",net0.n_7_3_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_5_zpos.txt",net0.n_7_3_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_5_zneg.txt",net0.n_7_3_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_6_local.txt",net0.n_7_3_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_6_xpos.txt",net0.n_7_3_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_6_xneg.txt",net0.n_7_3_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_6_ypos.txt",net0.n_7_3_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_6_yneg.txt",net0.n_7_3_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_6_zpos.txt",net0.n_7_3_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_6_zneg.txt",net0.n_7_3_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_6_xpos.txt",net0.n_7_3_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_6_xneg.txt",net0.n_7_3_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_6_ypos.txt",net0.n_7_3_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_6_yneg.txt",net0.n_7_3_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_6_zpos.txt",net0.n_7_3_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_6_zneg.txt",net0.n_7_3_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_6_xpos.txt",net0.n_7_3_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_6_xneg.txt",net0.n_7_3_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_6_ypos.txt",net0.n_7_3_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_6_yneg.txt",net0.n_7_3_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_6_zpos.txt",net0.n_7_3_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_6_zneg.txt",net0.n_7_3_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_7_local.txt",net0.n_7_3_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_7_xpos.txt",net0.n_7_3_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_7_xneg.txt",net0.n_7_3_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_7_ypos.txt",net0.n_7_3_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_7_yneg.txt",net0.n_7_3_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_7_zpos.txt",net0.n_7_3_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_3_7_zneg.txt",net0.n_7_3_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_7_xpos.txt",net0.n_7_3_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_7_xneg.txt",net0.n_7_3_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_7_ypos.txt",net0.n_7_3_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_7_yneg.txt",net0.n_7_3_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_7_zpos.txt",net0.n_7_3_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_3_7_zneg.txt",net0.n_7_3_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_7_xpos.txt",net0.n_7_3_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_7_xneg.txt",net0.n_7_3_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_7_ypos.txt",net0.n_7_3_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_7_yneg.txt",net0.n_7_3_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_7_zpos.txt",net0.n_7_3_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_3_7_zneg.txt",net0.n_7_3_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_0_local.txt",net0.n_7_4_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_0_xpos.txt",net0.n_7_4_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_0_xneg.txt",net0.n_7_4_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_0_ypos.txt",net0.n_7_4_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_0_yneg.txt",net0.n_7_4_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_0_zpos.txt",net0.n_7_4_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_0_zneg.txt",net0.n_7_4_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_0_xpos.txt",net0.n_7_4_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_0_xneg.txt",net0.n_7_4_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_0_ypos.txt",net0.n_7_4_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_0_yneg.txt",net0.n_7_4_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_0_zpos.txt",net0.n_7_4_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_0_zneg.txt",net0.n_7_4_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_0_xpos.txt",net0.n_7_4_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_0_xneg.txt",net0.n_7_4_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_0_ypos.txt",net0.n_7_4_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_0_yneg.txt",net0.n_7_4_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_0_zpos.txt",net0.n_7_4_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_0_zneg.txt",net0.n_7_4_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_1_local.txt",net0.n_7_4_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_1_xpos.txt",net0.n_7_4_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_1_xneg.txt",net0.n_7_4_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_1_ypos.txt",net0.n_7_4_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_1_yneg.txt",net0.n_7_4_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_1_zpos.txt",net0.n_7_4_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_1_zneg.txt",net0.n_7_4_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_1_xpos.txt",net0.n_7_4_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_1_xneg.txt",net0.n_7_4_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_1_ypos.txt",net0.n_7_4_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_1_yneg.txt",net0.n_7_4_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_1_zpos.txt",net0.n_7_4_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_1_zneg.txt",net0.n_7_4_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_1_xpos.txt",net0.n_7_4_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_1_xneg.txt",net0.n_7_4_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_1_ypos.txt",net0.n_7_4_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_1_yneg.txt",net0.n_7_4_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_1_zpos.txt",net0.n_7_4_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_1_zneg.txt",net0.n_7_4_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_2_local.txt",net0.n_7_4_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_2_xpos.txt",net0.n_7_4_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_2_xneg.txt",net0.n_7_4_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_2_ypos.txt",net0.n_7_4_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_2_yneg.txt",net0.n_7_4_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_2_zpos.txt",net0.n_7_4_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_2_zneg.txt",net0.n_7_4_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_2_xpos.txt",net0.n_7_4_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_2_xneg.txt",net0.n_7_4_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_2_ypos.txt",net0.n_7_4_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_2_yneg.txt",net0.n_7_4_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_2_zpos.txt",net0.n_7_4_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_2_zneg.txt",net0.n_7_4_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_2_xpos.txt",net0.n_7_4_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_2_xneg.txt",net0.n_7_4_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_2_ypos.txt",net0.n_7_4_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_2_yneg.txt",net0.n_7_4_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_2_zpos.txt",net0.n_7_4_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_2_zneg.txt",net0.n_7_4_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_3_local.txt",net0.n_7_4_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_3_xpos.txt",net0.n_7_4_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_3_xneg.txt",net0.n_7_4_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_3_ypos.txt",net0.n_7_4_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_3_yneg.txt",net0.n_7_4_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_3_zpos.txt",net0.n_7_4_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_3_zneg.txt",net0.n_7_4_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_3_xpos.txt",net0.n_7_4_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_3_xneg.txt",net0.n_7_4_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_3_ypos.txt",net0.n_7_4_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_3_yneg.txt",net0.n_7_4_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_3_zpos.txt",net0.n_7_4_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_3_zneg.txt",net0.n_7_4_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_3_xpos.txt",net0.n_7_4_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_3_xneg.txt",net0.n_7_4_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_3_ypos.txt",net0.n_7_4_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_3_yneg.txt",net0.n_7_4_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_3_zpos.txt",net0.n_7_4_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_3_zneg.txt",net0.n_7_4_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_4_local.txt",net0.n_7_4_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_4_xpos.txt",net0.n_7_4_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_4_xneg.txt",net0.n_7_4_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_4_ypos.txt",net0.n_7_4_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_4_yneg.txt",net0.n_7_4_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_4_zpos.txt",net0.n_7_4_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_4_zneg.txt",net0.n_7_4_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_4_xpos.txt",net0.n_7_4_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_4_xneg.txt",net0.n_7_4_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_4_ypos.txt",net0.n_7_4_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_4_yneg.txt",net0.n_7_4_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_4_zpos.txt",net0.n_7_4_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_4_zneg.txt",net0.n_7_4_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_4_xpos.txt",net0.n_7_4_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_4_xneg.txt",net0.n_7_4_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_4_ypos.txt",net0.n_7_4_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_4_yneg.txt",net0.n_7_4_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_4_zpos.txt",net0.n_7_4_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_4_zneg.txt",net0.n_7_4_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_5_local.txt",net0.n_7_4_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_5_xpos.txt",net0.n_7_4_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_5_xneg.txt",net0.n_7_4_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_5_ypos.txt",net0.n_7_4_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_5_yneg.txt",net0.n_7_4_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_5_zpos.txt",net0.n_7_4_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_5_zneg.txt",net0.n_7_4_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_5_xpos.txt",net0.n_7_4_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_5_xneg.txt",net0.n_7_4_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_5_ypos.txt",net0.n_7_4_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_5_yneg.txt",net0.n_7_4_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_5_zpos.txt",net0.n_7_4_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_5_zneg.txt",net0.n_7_4_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_5_xpos.txt",net0.n_7_4_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_5_xneg.txt",net0.n_7_4_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_5_ypos.txt",net0.n_7_4_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_5_yneg.txt",net0.n_7_4_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_5_zpos.txt",net0.n_7_4_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_5_zneg.txt",net0.n_7_4_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_6_local.txt",net0.n_7_4_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_6_xpos.txt",net0.n_7_4_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_6_xneg.txt",net0.n_7_4_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_6_ypos.txt",net0.n_7_4_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_6_yneg.txt",net0.n_7_4_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_6_zpos.txt",net0.n_7_4_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_6_zneg.txt",net0.n_7_4_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_6_xpos.txt",net0.n_7_4_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_6_xneg.txt",net0.n_7_4_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_6_ypos.txt",net0.n_7_4_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_6_yneg.txt",net0.n_7_4_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_6_zpos.txt",net0.n_7_4_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_6_zneg.txt",net0.n_7_4_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_6_xpos.txt",net0.n_7_4_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_6_xneg.txt",net0.n_7_4_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_6_ypos.txt",net0.n_7_4_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_6_yneg.txt",net0.n_7_4_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_6_zpos.txt",net0.n_7_4_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_6_zneg.txt",net0.n_7_4_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_7_local.txt",net0.n_7_4_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_7_xpos.txt",net0.n_7_4_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_7_xneg.txt",net0.n_7_4_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_7_ypos.txt",net0.n_7_4_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_7_yneg.txt",net0.n_7_4_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_7_zpos.txt",net0.n_7_4_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_4_7_zneg.txt",net0.n_7_4_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_7_xpos.txt",net0.n_7_4_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_7_xneg.txt",net0.n_7_4_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_7_ypos.txt",net0.n_7_4_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_7_yneg.txt",net0.n_7_4_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_7_zpos.txt",net0.n_7_4_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_4_7_zneg.txt",net0.n_7_4_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_7_xpos.txt",net0.n_7_4_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_7_xneg.txt",net0.n_7_4_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_7_ypos.txt",net0.n_7_4_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_7_yneg.txt",net0.n_7_4_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_7_zpos.txt",net0.n_7_4_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_4_7_zneg.txt",net0.n_7_4_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_0_local.txt",net0.n_7_5_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_0_xpos.txt",net0.n_7_5_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_0_xneg.txt",net0.n_7_5_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_0_ypos.txt",net0.n_7_5_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_0_yneg.txt",net0.n_7_5_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_0_zpos.txt",net0.n_7_5_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_0_zneg.txt",net0.n_7_5_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_0_xpos.txt",net0.n_7_5_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_0_xneg.txt",net0.n_7_5_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_0_ypos.txt",net0.n_7_5_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_0_yneg.txt",net0.n_7_5_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_0_zpos.txt",net0.n_7_5_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_0_zneg.txt",net0.n_7_5_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_0_xpos.txt",net0.n_7_5_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_0_xneg.txt",net0.n_7_5_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_0_ypos.txt",net0.n_7_5_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_0_yneg.txt",net0.n_7_5_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_0_zpos.txt",net0.n_7_5_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_0_zneg.txt",net0.n_7_5_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_1_local.txt",net0.n_7_5_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_1_xpos.txt",net0.n_7_5_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_1_xneg.txt",net0.n_7_5_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_1_ypos.txt",net0.n_7_5_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_1_yneg.txt",net0.n_7_5_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_1_zpos.txt",net0.n_7_5_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_1_zneg.txt",net0.n_7_5_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_1_xpos.txt",net0.n_7_5_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_1_xneg.txt",net0.n_7_5_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_1_ypos.txt",net0.n_7_5_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_1_yneg.txt",net0.n_7_5_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_1_zpos.txt",net0.n_7_5_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_1_zneg.txt",net0.n_7_5_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_1_xpos.txt",net0.n_7_5_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_1_xneg.txt",net0.n_7_5_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_1_ypos.txt",net0.n_7_5_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_1_yneg.txt",net0.n_7_5_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_1_zpos.txt",net0.n_7_5_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_1_zneg.txt",net0.n_7_5_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_2_local.txt",net0.n_7_5_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_2_xpos.txt",net0.n_7_5_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_2_xneg.txt",net0.n_7_5_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_2_ypos.txt",net0.n_7_5_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_2_yneg.txt",net0.n_7_5_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_2_zpos.txt",net0.n_7_5_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_2_zneg.txt",net0.n_7_5_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_2_xpos.txt",net0.n_7_5_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_2_xneg.txt",net0.n_7_5_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_2_ypos.txt",net0.n_7_5_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_2_yneg.txt",net0.n_7_5_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_2_zpos.txt",net0.n_7_5_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_2_zneg.txt",net0.n_7_5_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_2_xpos.txt",net0.n_7_5_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_2_xneg.txt",net0.n_7_5_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_2_ypos.txt",net0.n_7_5_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_2_yneg.txt",net0.n_7_5_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_2_zpos.txt",net0.n_7_5_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_2_zneg.txt",net0.n_7_5_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_3_local.txt",net0.n_7_5_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_3_xpos.txt",net0.n_7_5_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_3_xneg.txt",net0.n_7_5_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_3_ypos.txt",net0.n_7_5_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_3_yneg.txt",net0.n_7_5_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_3_zpos.txt",net0.n_7_5_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_3_zneg.txt",net0.n_7_5_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_3_xpos.txt",net0.n_7_5_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_3_xneg.txt",net0.n_7_5_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_3_ypos.txt",net0.n_7_5_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_3_yneg.txt",net0.n_7_5_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_3_zpos.txt",net0.n_7_5_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_3_zneg.txt",net0.n_7_5_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_3_xpos.txt",net0.n_7_5_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_3_xneg.txt",net0.n_7_5_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_3_ypos.txt",net0.n_7_5_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_3_yneg.txt",net0.n_7_5_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_3_zpos.txt",net0.n_7_5_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_3_zneg.txt",net0.n_7_5_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_4_local.txt",net0.n_7_5_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_4_xpos.txt",net0.n_7_5_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_4_xneg.txt",net0.n_7_5_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_4_ypos.txt",net0.n_7_5_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_4_yneg.txt",net0.n_7_5_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_4_zpos.txt",net0.n_7_5_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_4_zneg.txt",net0.n_7_5_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_4_xpos.txt",net0.n_7_5_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_4_xneg.txt",net0.n_7_5_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_4_ypos.txt",net0.n_7_5_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_4_yneg.txt",net0.n_7_5_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_4_zpos.txt",net0.n_7_5_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_4_zneg.txt",net0.n_7_5_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_4_xpos.txt",net0.n_7_5_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_4_xneg.txt",net0.n_7_5_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_4_ypos.txt",net0.n_7_5_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_4_yneg.txt",net0.n_7_5_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_4_zpos.txt",net0.n_7_5_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_4_zneg.txt",net0.n_7_5_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_5_local.txt",net0.n_7_5_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_5_xpos.txt",net0.n_7_5_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_5_xneg.txt",net0.n_7_5_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_5_ypos.txt",net0.n_7_5_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_5_yneg.txt",net0.n_7_5_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_5_zpos.txt",net0.n_7_5_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_5_zneg.txt",net0.n_7_5_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_5_xpos.txt",net0.n_7_5_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_5_xneg.txt",net0.n_7_5_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_5_ypos.txt",net0.n_7_5_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_5_yneg.txt",net0.n_7_5_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_5_zpos.txt",net0.n_7_5_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_5_zneg.txt",net0.n_7_5_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_5_xpos.txt",net0.n_7_5_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_5_xneg.txt",net0.n_7_5_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_5_ypos.txt",net0.n_7_5_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_5_yneg.txt",net0.n_7_5_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_5_zpos.txt",net0.n_7_5_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_5_zneg.txt",net0.n_7_5_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_6_local.txt",net0.n_7_5_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_6_xpos.txt",net0.n_7_5_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_6_xneg.txt",net0.n_7_5_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_6_ypos.txt",net0.n_7_5_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_6_yneg.txt",net0.n_7_5_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_6_zpos.txt",net0.n_7_5_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_6_zneg.txt",net0.n_7_5_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_6_xpos.txt",net0.n_7_5_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_6_xneg.txt",net0.n_7_5_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_6_ypos.txt",net0.n_7_5_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_6_yneg.txt",net0.n_7_5_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_6_zpos.txt",net0.n_7_5_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_6_zneg.txt",net0.n_7_5_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_6_xpos.txt",net0.n_7_5_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_6_xneg.txt",net0.n_7_5_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_6_ypos.txt",net0.n_7_5_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_6_yneg.txt",net0.n_7_5_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_6_zpos.txt",net0.n_7_5_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_6_zneg.txt",net0.n_7_5_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_7_local.txt",net0.n_7_5_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_7_xpos.txt",net0.n_7_5_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_7_xneg.txt",net0.n_7_5_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_7_ypos.txt",net0.n_7_5_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_7_yneg.txt",net0.n_7_5_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_7_zpos.txt",net0.n_7_5_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_5_7_zneg.txt",net0.n_7_5_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_7_xpos.txt",net0.n_7_5_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_7_xneg.txt",net0.n_7_5_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_7_ypos.txt",net0.n_7_5_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_7_yneg.txt",net0.n_7_5_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_7_zpos.txt",net0.n_7_5_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_5_7_zneg.txt",net0.n_7_5_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_7_xpos.txt",net0.n_7_5_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_7_xneg.txt",net0.n_7_5_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_7_ypos.txt",net0.n_7_5_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_7_yneg.txt",net0.n_7_5_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_7_zpos.txt",net0.n_7_5_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_5_7_zneg.txt",net0.n_7_5_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_0_local.txt",net0.n_7_6_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_0_xpos.txt",net0.n_7_6_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_0_xneg.txt",net0.n_7_6_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_0_ypos.txt",net0.n_7_6_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_0_yneg.txt",net0.n_7_6_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_0_zpos.txt",net0.n_7_6_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_0_zneg.txt",net0.n_7_6_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_0_xpos.txt",net0.n_7_6_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_0_xneg.txt",net0.n_7_6_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_0_ypos.txt",net0.n_7_6_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_0_yneg.txt",net0.n_7_6_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_0_zpos.txt",net0.n_7_6_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_0_zneg.txt",net0.n_7_6_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_0_xpos.txt",net0.n_7_6_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_0_xneg.txt",net0.n_7_6_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_0_ypos.txt",net0.n_7_6_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_0_yneg.txt",net0.n_7_6_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_0_zpos.txt",net0.n_7_6_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_0_zneg.txt",net0.n_7_6_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_1_local.txt",net0.n_7_6_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_1_xpos.txt",net0.n_7_6_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_1_xneg.txt",net0.n_7_6_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_1_ypos.txt",net0.n_7_6_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_1_yneg.txt",net0.n_7_6_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_1_zpos.txt",net0.n_7_6_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_1_zneg.txt",net0.n_7_6_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_1_xpos.txt",net0.n_7_6_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_1_xneg.txt",net0.n_7_6_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_1_ypos.txt",net0.n_7_6_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_1_yneg.txt",net0.n_7_6_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_1_zpos.txt",net0.n_7_6_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_1_zneg.txt",net0.n_7_6_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_1_xpos.txt",net0.n_7_6_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_1_xneg.txt",net0.n_7_6_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_1_ypos.txt",net0.n_7_6_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_1_yneg.txt",net0.n_7_6_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_1_zpos.txt",net0.n_7_6_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_1_zneg.txt",net0.n_7_6_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_2_local.txt",net0.n_7_6_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_2_xpos.txt",net0.n_7_6_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_2_xneg.txt",net0.n_7_6_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_2_ypos.txt",net0.n_7_6_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_2_yneg.txt",net0.n_7_6_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_2_zpos.txt",net0.n_7_6_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_2_zneg.txt",net0.n_7_6_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_2_xpos.txt",net0.n_7_6_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_2_xneg.txt",net0.n_7_6_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_2_ypos.txt",net0.n_7_6_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_2_yneg.txt",net0.n_7_6_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_2_zpos.txt",net0.n_7_6_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_2_zneg.txt",net0.n_7_6_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_2_xpos.txt",net0.n_7_6_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_2_xneg.txt",net0.n_7_6_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_2_ypos.txt",net0.n_7_6_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_2_yneg.txt",net0.n_7_6_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_2_zpos.txt",net0.n_7_6_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_2_zneg.txt",net0.n_7_6_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_3_local.txt",net0.n_7_6_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_3_xpos.txt",net0.n_7_6_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_3_xneg.txt",net0.n_7_6_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_3_ypos.txt",net0.n_7_6_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_3_yneg.txt",net0.n_7_6_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_3_zpos.txt",net0.n_7_6_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_3_zneg.txt",net0.n_7_6_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_3_xpos.txt",net0.n_7_6_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_3_xneg.txt",net0.n_7_6_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_3_ypos.txt",net0.n_7_6_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_3_yneg.txt",net0.n_7_6_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_3_zpos.txt",net0.n_7_6_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_3_zneg.txt",net0.n_7_6_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_3_xpos.txt",net0.n_7_6_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_3_xneg.txt",net0.n_7_6_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_3_ypos.txt",net0.n_7_6_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_3_yneg.txt",net0.n_7_6_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_3_zpos.txt",net0.n_7_6_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_3_zneg.txt",net0.n_7_6_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_4_local.txt",net0.n_7_6_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_4_xpos.txt",net0.n_7_6_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_4_xneg.txt",net0.n_7_6_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_4_ypos.txt",net0.n_7_6_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_4_yneg.txt",net0.n_7_6_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_4_zpos.txt",net0.n_7_6_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_4_zneg.txt",net0.n_7_6_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_4_xpos.txt",net0.n_7_6_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_4_xneg.txt",net0.n_7_6_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_4_ypos.txt",net0.n_7_6_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_4_yneg.txt",net0.n_7_6_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_4_zpos.txt",net0.n_7_6_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_4_zneg.txt",net0.n_7_6_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_4_xpos.txt",net0.n_7_6_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_4_xneg.txt",net0.n_7_6_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_4_ypos.txt",net0.n_7_6_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_4_yneg.txt",net0.n_7_6_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_4_zpos.txt",net0.n_7_6_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_4_zneg.txt",net0.n_7_6_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_5_local.txt",net0.n_7_6_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_5_xpos.txt",net0.n_7_6_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_5_xneg.txt",net0.n_7_6_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_5_ypos.txt",net0.n_7_6_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_5_yneg.txt",net0.n_7_6_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_5_zpos.txt",net0.n_7_6_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_5_zneg.txt",net0.n_7_6_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_5_xpos.txt",net0.n_7_6_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_5_xneg.txt",net0.n_7_6_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_5_ypos.txt",net0.n_7_6_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_5_yneg.txt",net0.n_7_6_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_5_zpos.txt",net0.n_7_6_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_5_zneg.txt",net0.n_7_6_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_5_xpos.txt",net0.n_7_6_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_5_xneg.txt",net0.n_7_6_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_5_ypos.txt",net0.n_7_6_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_5_yneg.txt",net0.n_7_6_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_5_zpos.txt",net0.n_7_6_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_5_zneg.txt",net0.n_7_6_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_6_local.txt",net0.n_7_6_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_6_xpos.txt",net0.n_7_6_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_6_xneg.txt",net0.n_7_6_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_6_ypos.txt",net0.n_7_6_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_6_yneg.txt",net0.n_7_6_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_6_zpos.txt",net0.n_7_6_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_6_zneg.txt",net0.n_7_6_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_6_xpos.txt",net0.n_7_6_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_6_xneg.txt",net0.n_7_6_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_6_ypos.txt",net0.n_7_6_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_6_yneg.txt",net0.n_7_6_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_6_zpos.txt",net0.n_7_6_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_6_zneg.txt",net0.n_7_6_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_6_xpos.txt",net0.n_7_6_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_6_xneg.txt",net0.n_7_6_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_6_ypos.txt",net0.n_7_6_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_6_yneg.txt",net0.n_7_6_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_6_zpos.txt",net0.n_7_6_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_6_zneg.txt",net0.n_7_6_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_7_local.txt",net0.n_7_6_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_7_xpos.txt",net0.n_7_6_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_7_xneg.txt",net0.n_7_6_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_7_ypos.txt",net0.n_7_6_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_7_yneg.txt",net0.n_7_6_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_7_zpos.txt",net0.n_7_6_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_6_7_zneg.txt",net0.n_7_6_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_7_xpos.txt",net0.n_7_6_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_7_xneg.txt",net0.n_7_6_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_7_ypos.txt",net0.n_7_6_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_7_yneg.txt",net0.n_7_6_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_7_zpos.txt",net0.n_7_6_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_6_7_zneg.txt",net0.n_7_6_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_7_xpos.txt",net0.n_7_6_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_7_xneg.txt",net0.n_7_6_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_7_ypos.txt",net0.n_7_6_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_7_yneg.txt",net0.n_7_6_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_7_zpos.txt",net0.n_7_6_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_6_7_zneg.txt",net0.n_7_6_7.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_0_local.txt",net0.n_7_7_0.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_0_xpos.txt",net0.n_7_7_0.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_0_xneg.txt",net0.n_7_7_0.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_0_ypos.txt",net0.n_7_7_0.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_0_yneg.txt",net0.n_7_7_0.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_0_zpos.txt",net0.n_7_7_0.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_0_zneg.txt",net0.n_7_7_0.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_0_xpos.txt",net0.n_7_7_0.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_0_xneg.txt",net0.n_7_7_0.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_0_ypos.txt",net0.n_7_7_0.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_0_yneg.txt",net0.n_7_7_0.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_0_zpos.txt",net0.n_7_7_0.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_0_zneg.txt",net0.n_7_7_0.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_0_xpos.txt",net0.n_7_7_0.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_0_xneg.txt",net0.n_7_7_0.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_0_ypos.txt",net0.n_7_7_0.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_0_yneg.txt",net0.n_7_7_0.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_0_zpos.txt",net0.n_7_7_0.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_0_zneg.txt",net0.n_7_7_0.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_1_local.txt",net0.n_7_7_1.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_1_xpos.txt",net0.n_7_7_1.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_1_xneg.txt",net0.n_7_7_1.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_1_ypos.txt",net0.n_7_7_1.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_1_yneg.txt",net0.n_7_7_1.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_1_zpos.txt",net0.n_7_7_1.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_1_zneg.txt",net0.n_7_7_1.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_1_xpos.txt",net0.n_7_7_1.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_1_xneg.txt",net0.n_7_7_1.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_1_ypos.txt",net0.n_7_7_1.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_1_yneg.txt",net0.n_7_7_1.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_1_zpos.txt",net0.n_7_7_1.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_1_zneg.txt",net0.n_7_7_1.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_1_xpos.txt",net0.n_7_7_1.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_1_xneg.txt",net0.n_7_7_1.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_1_ypos.txt",net0.n_7_7_1.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_1_yneg.txt",net0.n_7_7_1.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_1_zpos.txt",net0.n_7_7_1.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_1_zneg.txt",net0.n_7_7_1.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_2_local.txt",net0.n_7_7_2.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_2_xpos.txt",net0.n_7_7_2.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_2_xneg.txt",net0.n_7_7_2.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_2_ypos.txt",net0.n_7_7_2.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_2_yneg.txt",net0.n_7_7_2.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_2_zpos.txt",net0.n_7_7_2.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_2_zneg.txt",net0.n_7_7_2.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_2_xpos.txt",net0.n_7_7_2.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_2_xneg.txt",net0.n_7_7_2.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_2_ypos.txt",net0.n_7_7_2.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_2_yneg.txt",net0.n_7_7_2.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_2_zpos.txt",net0.n_7_7_2.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_2_zneg.txt",net0.n_7_7_2.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_2_xpos.txt",net0.n_7_7_2.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_2_xneg.txt",net0.n_7_7_2.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_2_ypos.txt",net0.n_7_7_2.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_2_yneg.txt",net0.n_7_7_2.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_2_zpos.txt",net0.n_7_7_2.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_2_zneg.txt",net0.n_7_7_2.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_3_local.txt",net0.n_7_7_3.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_3_xpos.txt",net0.n_7_7_3.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_3_xneg.txt",net0.n_7_7_3.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_3_ypos.txt",net0.n_7_7_3.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_3_yneg.txt",net0.n_7_7_3.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_3_zpos.txt",net0.n_7_7_3.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_3_zneg.txt",net0.n_7_7_3.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_3_xpos.txt",net0.n_7_7_3.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_3_xneg.txt",net0.n_7_7_3.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_3_ypos.txt",net0.n_7_7_3.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_3_yneg.txt",net0.n_7_7_3.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_3_zpos.txt",net0.n_7_7_3.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_3_zneg.txt",net0.n_7_7_3.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_3_xpos.txt",net0.n_7_7_3.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_3_xneg.txt",net0.n_7_7_3.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_3_ypos.txt",net0.n_7_7_3.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_3_yneg.txt",net0.n_7_7_3.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_3_zpos.txt",net0.n_7_7_3.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_3_zneg.txt",net0.n_7_7_3.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_4_local.txt",net0.n_7_7_4.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_4_xpos.txt",net0.n_7_7_4.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_4_xneg.txt",net0.n_7_7_4.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_4_ypos.txt",net0.n_7_7_4.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_4_yneg.txt",net0.n_7_7_4.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_4_zpos.txt",net0.n_7_7_4.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_4_zneg.txt",net0.n_7_7_4.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_4_xpos.txt",net0.n_7_7_4.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_4_xneg.txt",net0.n_7_7_4.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_4_ypos.txt",net0.n_7_7_4.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_4_yneg.txt",net0.n_7_7_4.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_4_zpos.txt",net0.n_7_7_4.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_4_zneg.txt",net0.n_7_7_4.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_4_xpos.txt",net0.n_7_7_4.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_4_xneg.txt",net0.n_7_7_4.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_4_ypos.txt",net0.n_7_7_4.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_4_yneg.txt",net0.n_7_7_4.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_4_zpos.txt",net0.n_7_7_4.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_4_zneg.txt",net0.n_7_7_4.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_5_local.txt",net0.n_7_7_5.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_5_xpos.txt",net0.n_7_7_5.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_5_xneg.txt",net0.n_7_7_5.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_5_ypos.txt",net0.n_7_7_5.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_5_yneg.txt",net0.n_7_7_5.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_5_zpos.txt",net0.n_7_7_5.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_5_zneg.txt",net0.n_7_7_5.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_5_xpos.txt",net0.n_7_7_5.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_5_xneg.txt",net0.n_7_7_5.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_5_ypos.txt",net0.n_7_7_5.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_5_yneg.txt",net0.n_7_7_5.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_5_zpos.txt",net0.n_7_7_5.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_5_zneg.txt",net0.n_7_7_5.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_5_xpos.txt",net0.n_7_7_5.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_5_xneg.txt",net0.n_7_7_5.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_5_ypos.txt",net0.n_7_7_5.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_5_yneg.txt",net0.n_7_7_5.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_5_zpos.txt",net0.n_7_7_5.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_5_zneg.txt",net0.n_7_7_5.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_6_local.txt",net0.n_7_7_6.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_6_xpos.txt",net0.n_7_7_6.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_6_xneg.txt",net0.n_7_7_6.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_6_ypos.txt",net0.n_7_7_6.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_6_yneg.txt",net0.n_7_7_6.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_6_zpos.txt",net0.n_7_7_6.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_6_zneg.txt",net0.n_7_7_6.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_6_xpos.txt",net0.n_7_7_6.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_6_xneg.txt",net0.n_7_7_6.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_6_ypos.txt",net0.n_7_7_6.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_6_yneg.txt",net0.n_7_7_6.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_6_zpos.txt",net0.n_7_7_6.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_6_zneg.txt",net0.n_7_7_6.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_6_xpos.txt",net0.n_7_7_6.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_6_xneg.txt",net0.n_7_7_6.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_6_ypos.txt",net0.n_7_7_6.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_6_yneg.txt",net0.n_7_7_6.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_6_zpos.txt",net0.n_7_7_6.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_6_zneg.txt",net0.n_7_7_6.switch_inst.ZNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_7_local.txt",net0.n_7_7_7.local_unit_inst.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_7_xpos.txt",net0.n_7_7_7.switch_inst.XPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_7_xneg.txt",net0.n_7_7_7.switch_inst.XNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_7_ypos.txt",net0.n_7_7_7.switch_inst.YPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_7_yneg.txt",net0.n_7_7_7.switch_inst.YNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_7_zpos.txt",net0.n_7_7_7.switch_inst.ZPOS.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/routing_tables/routing_table_7_7_7_zneg.txt",net0.n_7_7_7.switch_inst.ZNEG.routing_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_7_xpos.txt",net0.n_7_7_7.switch_inst.XPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_7_xneg.txt",net0.n_7_7_7.switch_inst.XNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_7_ypos.txt",net0.n_7_7_7.switch_inst.YPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_7_yneg.txt",net0.n_7_7_7.switch_inst.YNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_7_zpos.txt",net0.n_7_7_7.switch_inst.ZPOS.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/multicast_tables/multicast_table_7_7_7_zneg.txt",net0.n_7_7_7.switch_inst.ZNEG.multicast_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_7_xpos.txt",net0.n_7_7_7.switch_inst.XPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_7_xneg.txt",net0.n_7_7_7.switch_inst.XNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_7_ypos.txt",net0.n_7_7_7.switch_inst.YPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_7_yneg.txt",net0.n_7_7_7.switch_inst.YNEG.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_7_zpos.txt",net0.n_7_7_7.switch_inst.ZPOS.reduction_table);
	initial $readmemh("C:/Users/Jiayi/Documents/GitHub/MD_reduction/tables/reduction_tables/reduction_table_7_7_7_zneg.txt",net0.n_7_7_7.switch_inst.ZNEG.reduction_table);
	initial begin
		clk=0;
		rst=1;

		#100 rst=0;
	end
endmodule
